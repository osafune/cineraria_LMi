��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�=�}A1��=1�<��xr7�n�?��;�MHc ��c��Ɨc�ɍ|�w1�ag�j�J�gDBʚ��n�N���a�� Zs��Gb��'�[����_��.#�2��*���|�PNž�0t��'�֩�X~!���i0��A��-�xI'O:1�T���v��W�r�� u���ڍ3�����G����Lֿ�^PQě��zg�nJ����*��EV�I�����u�杇�e,[��l��9Љ�`u6���4�
R�ox�uT\)F�^a�¦/��`ɁK�<��]Ñ�tt�GGe��[�]GO���Ŵ_Kb��f�Ok�i�(���\�,��br;ғD����1�Q������$7�N�����S?L��:�sJ}��%oy��������3�ڴ`��?�le�9��<m�P�y�!�!��sN�E��k�+h�602y�n�AtW�����V��N�"{�042'3����L��l�d���E�3�����Li�&3�����o�����Kk��:h�A�,:qoB�qU�g/�_a1hl���vo�$v����3��4�?-N[����w ���nG2ڻfod�<m�)�������h�x���n.��q��R��^�w5��76�� �8�m<�.U�@�:���i���jH��Ex�Ю���N����.�5p�V�l^�������Ft=֧@{�k;Ee�y�դ��K��Y%��b�ĸA;�QC:��������F��c�A��д�~I��O�,kL�S���q�eH�R����܅�g�2ۺW�M���?�!���;��b��\v|�d����^^�Ȱ�[��r;�e�WN��b���t�w���KĬ��O�y���-�gYդ����m�3�Fbպ����u�@�TE����Ȳ��#���I�>Dں�GgQ�`(��	� `������H�p���X��X��i9p�s��jCLa�'rg�_���ZǪ@��fͨ-�����Ia�a�i[�73����$��.�5��Y�׼2��KÒ�y����$��\�M�/�s��s��4�37��Q�%z�O;h�T_cm4Ӈ��*x��}SaV��`Z�C�%mdt��\��)�}�S%�5�Dh��%>]�H�*�<��_B�� ���]��O�J����[D�B�}�F�gq�-��tb�8�~���*��r�q�r��J/���x�*�ܗ>�����T��ƿ3�b�a;��O�*j����*F�� RO4�p��Y7+��1��q2D�`#E2�^I��U��É�4�*�S�{9��zykhA-�ɛՀ=�����.�q�3�`�x2�6��ln�C޳�!�\-I#kP��][
7l��'��R�I~�Ǌͅ?:jn܉���|�(q����{y�R��(@M��Tj��N�6���Q���E�`�w��i��][���� �IXǀfg�v��}�Rt#��R�x���&��<a�s v��������%H�ځ�48M�/�_]M���Ɣ��U�y7�B��H8h��D|P9K�1�3{�W����N�pؾa�@�
���}��U��R:�!�*yO��l�K�������.ؠ�8�A�zӖK���Gws� D �mF�,1_���S^J�/��{�xT�q���y�Y�Q���E��H2񇼥;����_�';�?���{�vR@J�EF�����`�V��nͫX��`<x[B
�	Oϱ�<y;�`ѻ�IOÅ\��Yf�V~SC8����#���Te�m7�n�,s��,���CׯZ$�Mg��/l�=l���s�+R���bʃ�	�����x��i|F�,5��n nK�e���k"��Q�0[�+��/�7v�Z�5�Re��S���7�^h�g�8�G2��NKZ�Xٲ�c�J.�Gb2SQdg�I@0n=P�i�{}�pK�H��n�M6��y86����[)?�.UR�M:���	Y��A�r2��r��{��_��=�Эa��sM�E��\{C)���w<I#�Q��Q�8�DS��(!]�F긹
{����k�׭)�AIw�[������Y�^����g�eP���)W��~�[�D6j��w��:}�}9 �D�'�,�E�.��9�� ��6	��%2:G`��t�X�LE�gd�U؆ә3�cJ��g!�-'���<���0<K���Mg�BH��7��_��1�/��W[6A���1��}�)��m�G!�^D}��MW��\�N5��7���?�t ��H?V������`&"?/ͯ�v�����r˕L��u���,�nX���b[N���x���Z��Fͥ��f�a�u��h��c��T؝�L�lM�4�!IuW�˽� �/t���3qH��d�cVL+����ֈ�{'=b0if���Dٿ���s��kQ$p��N��#K�aLiC+@��
��;>S1&���ݜ�O;�o�u$i����6�Wr	~�Q0.���Ԝ�E��a��K���:-Foz�z%��6��Ɋ9����!i�6�:$����7
k~�i3�S7@�g��5l�9�����,>����WUl#�ǹ��m��GZ4|�LM�0�qx}�٤rY*Ǆ���0� #���Wu���yˡ�ۡ���ϥ�5�P#>�����c�s;]�<�+<�2���#ec)�\�ʒ}��D�.ye���J:��Ĉ&���Yj����DQɨ�gE\������.�
����[FPt�>a�_� ?��-Mk��fc(T*UĲD$�OɮE�B�D����zq^�T}�����n�b�#�2��\�M�vF�.���.[��<^���dNu�K#6�	~q�Yj�9���Pyq�h}�FY�W��I�������J3d��%�W�S������R[K['`8)sm0�I�Wi��~(QPmCw`�����@���2��݈�o��ĥ�8^+�֖wh��`���%?G��+K�����7��daLo|>���ݻܨ�੫��Z�PCN��}dO� �9,Z�_��ʹT��<�# /�1tpjߌ�bU�7�<�C<F/i�q+eqw��U#|ibt�+�X�7O� ���Ȃ�	����s%7�ŀ��!��{���[웤P�4Ax6щJ�Z�\�p�FS8��dn����|@XWLW�Ht�O�Ա|x�퓦�d��sB%A���'���S:$��U�&θ1HW�Q�/�����%�l��Ջ�OjSH̵UKA����4�7�R�D灯��������Hǩ
���m|]/�� (7ݻ���ǦϹP2���r�O@H�/P+r�����L�<G䦮�XF���h��Q�G�Jkko�%������Fv�̊).hxz�d/���\�+�*��L�>N�(�QA�m�V �>f��c|5�,�y��QȟYԻL�c�$�.���Z��d��P�C���n��w���QXO��@��.	B�^�ae�;�1ذ�<D��_8N�:b����Q!|��IQ5561l��d���=g�>�gSxgew�e�Y��c~�'��?�N�gȕ��
X�f�l��[y1��-���������3��g#;7
,�g����p9*$�o%��~��s��Vŋ�ϩ/?fh��򊀜�n�B��������S��8�*�<~%�ۆ���[1�{'JoH�v����K�Z���ɲ�)� IƏ�sB����"oI]qZ���P?���6��#�մ�ǃ��b|��L��KaP'�;�F�d�}���_F��yO��Jl��4�r�J�~F��w&���Q�qz�.�'���6�'�J��=�^�]�%6�2�(����E�#�t�"���E��JZ4.�ę����[����m�(�H.���V��?���ӱ��(�b,6�RD�O�$x>�0)���T5��f�4��W�=o��}�w�t,�0�r<=��������i����P0�7�1��LD���f �۔s�9T�Ֆ�a�D�5��O�峐��#=��1�M�Jbv�?;��-j��ø�O���f5�nE{�6s�L�j�I5%�,w��g�s�}�^��P"f�A�O��c�P+��z���u�Aj]�؆�19,L��m�v���Ț=~��R$����IhW;M��>I�����I����pK���A x�	x��I̩���Ĝ�Ul^�4kV8���)�P����.��V�1,P!��Z%B��Ы��G�N;���cn�h����.R���_�oʵm�h��V�MP���Z7��G,�#�K�Y9-N�yS�`:A���->LkƀK���}�XݑX�prI�=I�C4�h�0�Л�o��`/V�Q����Y3�+�~�*ۿ	T�
���c"��ՠ�y2K��9@5ꐮh���E�M6@A ���=X���}�2�)���Zʣb��&��+8��vb &���_��p0�I�v��R9��H�C=����������S^4�Yp��=I(36w��%�A?��S�%|��x�mL`�a���D���p�7,�(W��z�=�D#-&w֨��<��`�B
gѭ)�$���I)���BPv��ɊCg(��u�؎a*�x]R&rw���4l�tQ��x@������H��d[��aO��̭���K쉶�H�2�<]�W)�
�����۬gdpg�=�1��4L���;�QUp�[��ݤ�o�� ��a4�7��o���~��Ϋ���K/�H�xǮz;te�(8���\�)U�8���P��N���+D�`�3	&$��GO�{[u� �d�ו}��B-���yr�=�ׅ�"}2?�Di�k�΂hO�r}/��Rwk6���n���9w���ZO�����p��ȭY�vɗxrq���R�W�t���M�^�Q|B��W����H�����5��T��&>�d|4}%T!���J�T-���Pwo�x$��VIa��d��4���#��{.��t�Ч�V��y��@�  �����tz�����6��\��+.� D!�\���#�G�g�,%�+�s������Ə����{�٠p��暜�WuMO��Q�8�8�ۭ�� � zt��"��ݔ��a!��%���ҩ��ȬE&Ҁ�[��>�~��]�pL�M1x憁��fo�AY��0�r�����C�d%�mX���[\��\�I�좒O��2 0�8s�,@
݈��h{�v<�cK�8HKg �YAZ�	I�P��U�c����ߐM����`�˿t�)$��4�������*���w#��Wx��_ul�[%3��i	��4�9r��S: G�B���a�6�g�ۚ\����ȫ����1d������'��P��X,]Y���o�� êd���P�Ex�4��pW�o뭳#Z�=/ho#�X����,��W �/Gׁ�!����6f�9A��u�AА�"]��J���n��X����p|�L+��Cg��#�����=��v ?��u�����yhT�0�7������f�E&�#	$;r�Bp�1��3��9�+�g�m�$(PRA�
��±���
���ł�����e�;d��K8��&�E����Y���I���h�+ۂ�dDґ����~Y����q�J�s\�=�	�Pd[Մ��]�%��3�l�!�Q_+�t&���g�x1��	у�}A���3�y\���5�A��?��|L�U��Dx0c���
����d��J��Q�i��3қF�x�����#��	����B<�W/E�|�_By�Y5�㦊�D��Pgi Ʋ������L ��P׽/��g>�5��Z�5�;�,��R��]fm�_�cc|�Ҙ�k�n5�ՀTċ��h��9&z��;��T�*��	�}Q@!-��-���yt��B�1���6��^7�Cq�A���7��ʸ�������@�v�dp�[V������wE�<Ѱ�Wb"���A��vZ�� ���㍋�s��
�!d�̑҃�l'�T&VG�R5DE`upHУ����z��5��2��a8�{ˀ�c�k��Nn������cȮ+���EL$��#C&�P�d9v�� 0����R�L�H��U{���X��d\$�م�晨O������w뜌�| Ba�����?�l~x=��/�Abx�#�?-:�	3��_���捡�tRiv�����$��}>�׊��`Y��#�U�N�zD$���F�)�|�&�(f�&�d��~� Z�k�׬{C+fmo�B]��ܲ�cK�^�e�o@kA��Xѻ��5�2�1P=u��͈~�Uޘ:B<�|��uLCPH��CUyrZ�F�"����/�E�p�D���ƂWK���K&��9t!(��Q�揙���U��yF�.(�v�=����);��R��|��D�en�燇ƞ���BGD�#��U�L�ߛ�>auQ�����]��~]<"ǹ�("��׳5Gv���ee}����*�;
�ئ��a
v��ۭ/�q��,�c���W�t���������6`�/by?>��[��T�{�����T�z�� *��֚������~
�1+j���NS{��<�s��#��5��Q��tӾ�|v�� K/�MGh�߄_�:$���?��� nG@#bva�Y�r΀�^�|eXΣ
�\_Y՟9�8g?hژ���Ʒ����նKY��c=���3�-Lo=���Zq�c�Ƀjss��7 �WbD=��zʴ�Ӗ(��À����F���@G��� ��AU��s�C�<�L�.��d���Oxt ��.��8��{hI�(�������-,��1)������6����L>���V��u!L������_�������1G\Wo��RV#�
N�w&�`��9�z�!�*7-��� ��4�~�iN������&�4���A�$����Pa:z8}�p���A�-��h����2q���сb-����3Lib;�֤�B��-A�����V O��p���@��v�N�3	�BZ;�%5�p������O��x����~�{�|�����~��xi�
���a�Wt:	e�U8)0�m��A]��Q�^�i�<��>-q�Kns�*�L���l�%v T����'��/L�#��εoS������H��rf2/Q ��ff�J#΅�M�wY�@+����&B�X^e�hZ����}�󥼁�"J;e�o4y	��>��0�����#���
���$EpVz����b�M����Z!6_�t���B��v�+F��ع-�7�z_E�K|/��y��洡����v��+Z����r.�` T%����n�d^Y�Ŝ���q0�ؕN��t��|��4�n]<{��=�����˗p�D�a�P=lF3��݄4;:���5�6�^]�xODˇ������Ir������-Y�lB��"5�93�V��]�3�m(��FU��H�^߄7Aj$|�O�c�2�n
������u8� ,����������G���5�<����w�k��1�m��E�	ˀ�2�o��n��ūT���H/�5\-1jݧ%�ydE�O�_D� ���X��7�>������)N8� �/�	nf �A���
��~�O�v�]3�I�4�[�g���gb�q6n׆pD�sJ�&�*n`*�_z��`/?�<�����]4I����
�*� �~Mv�}��*IW�v�7;��XN���G8��X�K(�@�OF��֘��e�1�;nZg���?׎)�>%\���u5em���'1�3]��9Ԛ>��p�>�Iڰ3�����g%RO*�>�C ����O��l��Ku�y�� ����#�}��g�fW�����ͥ��D���	t���.�,�'��Տ����s'eADh�Ɩ��}��h�eO�ow^�F�Զމ���ߪ{D0���v��$�~I�h՝��T�!��?DR�n���>R^��L�[(3����s�v� �ЛZ�A0B�d��Z�,����/�{s�/�ce��H�~:�Ȋ�P���i�9�)dH(���(V�,��k����t�;��F��#�)#�IŵS 2s��S�w拭J�	 � |�Q������� ʹ�&�U�l�6�M���

�d�f"���S�x��E}����۱V8��)�~0�?���+�G۩΃���i�5O#4a-mB��Q�ϖ��'�E4L��8�~O5��1 +��8���8���p�iN�a�pY����V��69�f;��H�Ґ-<�o𣬈���'-p�px����m3KˆX�B�P]�\	�o(�}p(��PM��$�����,A�@,yk:d[$p����ߋ���uC�8�i��Y]#+Q�E��H��O��i����p_�g3��&[7��Ĭ�x�d�Y�x�:�cI�$�(���#�-�����p�w�BJ͋ږ�uz �����t{��6t��l���*e��'_������`c��C�Z���'!"���8��s��w��f~@���.�x�����A��<�css�2�C�E���GY�2����,�sW=V���0�J���~Z�(�%�0�`J.����@��`�M�C�2Z�!�|xG�r`3ԙW����9Q�ub�ਰ�u;��q�ն���Ωؐ][9p�v�����E����Y^#���G�|IְR��</�jm��j�*�뾳)ñ�+�}L�����MJ�`��l�b�����lG�Z����<���*�(�+Z���|�Q47䨸&&�&�Y��=������*��w;�3�8͇l 9t��<��<hïƧ洽�*e��gqg������j�Ly,���EJ��D��Q��e�4p��S�DE�&i��a�8�V��u_��x P@�t#7*�l��=���F�̌$r����MMC�&c��a�$�����ߩ�B����݆��r�w�6��K0�Y��>�F��*��	�8�~qB�-7���v���%�&�!%䊗8�H�W=8����	�t�q�'�D(����9�xCy YР��z	F
�"Q�^��*w9;^��Ű����_�>l��^��=��~9�e�-"r�P�|%j��
6�`Ƃ�����싈�/�<1�����[�ƀ��(g�)�%;j����<����X!��]^��I#�QIN�����Oh;�v�s����g��'�c� ��XE�ik\�ͣ�2G�Y(���ʙ(H�F����K����)*1!�\��4�6�*;0i�s`��{A�`M8���B��|��3&��Zպ_�wC��1��������$K ��h��������ұ�E��m�� �0����H�௭��)�:��Jh�/�i�q�x�yz�f���߸|��<TT�	�e�Z�����g����9+�/ڭ�BA8�/T�%g���~m��%����a��HP�]E�c@�R#�o�ͭrդ�%�~��!Q^��l3����.���V���/��K9P ��I�,��
L�Uc&|���7WT���/h0�ef#������yd�'$�7c�0��(���+����3�W}��*���]T�ݙ1�?Yy��6�c�ߖ[/½˞�����NA1\�Sж��Wk��	�o����tZ�ah�A�K��Mm�]�o�:��ҷh���nzB̏�BVsP�U��X�VVi��߈�q�L�LXp?|N��M>͞��ԫ�PIP��Y����Pa4�z�1*�.��f�����"�U��|fYz��� ?<8V�eM�i��QG_?���v�Hn�j�&�������XhPlV�8Z��W}��XSt�-��z�Hq=P��C,�m���-��pI%4Q���2�޹���qXc��sv�*p�/Zy��
6�[�D�9Y3C¿��q�x�v41+#ڸ�F��6�wi�T�Y^x&>Y�g��̱
ا"Л�n'��:yU���WO��u.�F֯������eeN�ab�Zx�$�$g�m�Nu|�߾��3�i|�(�ƞ����}>�d8wWe���m+�ұ<ʼ�5�����%ji����W�h���'�6������;5r��FL�81P�g�RH(]�_V�+!9k���dhc#VxwP��H�D#`X]�t��q�u�'��vP���F��(�1Ğ�?�MQ�uO�3ViMvm��^
_rJ&獸ɱ�wK\L	vUV�W�m��_� ae\/��a���Uz��{�ގ�0�/=����~��8�oY�>�!=��xMU�2��<%��9���	�O@����ţ�W���J޹A����͜�v:s�����g�R�w==v��|Ié�@5���Ϙ5�QP��z�\ ���<�x��0���F��tw�S�_>� iwE�@��O���� �5w�p?����~� ��e���9���쿨�f1����SQʩX�> y���[���Xr��[�Ņ�C�ܾ>��Y� ������F��<��l��g@���� ��֡Z��������i�)�5�b6zy�-�m[�]tOI���k�E|��P����^��]��<c�I���FSI���@���L�JZ�I+8}X��U+W.��snzP��� ��u��2��}�T�m`^�p��DSQ|�Oɐj���F4�w��bġ��US�}�*N�}�8q���Z�ھ�P� ߛ�n��3��eF�����0��-�B Aʧ�bVQ4�UF�������Sm����׀U�bk��;^�p���7�R^O�(����0�$�5k2��P�$z�?I	�c����x7ρb���i!�"��x~h7]Sģ�-�~�[#�o��,T�	���܀�Ob������(%UmO��O��������{�;-�JJɈ�X鑅Y۔��1�n���Q
Wh�ޱ{3n'�_���� gJ�>�
�tG�����_-�Ľ�h�͒*��p˄��3���!D<��A���L��%:�]\�nZ��!���I�#���Ąw��u�D?+Ly�ۼ$`sk��;\��&d�٩"��-�"RO�6�;�!�u��ID���N�D�_Sdc"�b`]��L�$\)��ʧ�]'���<h��d SzE߿��8IY`��e
P:cͺl�67����M�+�^ks%anR�ڹs��H�,p!ψ�!X	к��̘��g�Ĵpu%��%WK�}=4H5_��Uu��߸�C�Oj%�դ���8Sye��5�T]Am.�f�P����xBP)|�+e�"�ؿƥ5�j�^u����Dć���P�=J����>$#6��������a/�px7�l�*
�z�_I;F�E⻴�?�3q։@�t��s�;�`h;� �����\~B�â��b�b:�k�#�9A#����Ĥ�6�v\�?����l��ԳB6֪6����R�� �𧦛�y{�Qg#��#Z��m�9Q'\�K7�sʜ3}��-JU��p*�QI��#�p��2<�#����;�LߴЇ4��,��t�<�'สE��O"s]�"(����u�R��*V,�U����NZċ8�%<�s��u�3@���~*h��V�@Ou��oj?��#���+���7���}�S�7�_�P,Ze:A7�� R��e��3L8IvT�h��-Aע�v���M��r*z����~�{��ԅ��X�^,M-�rm��Y�sW</�X����Z}��-��+G��s5���F�,Fy�5��wdIu_��������S��"�H��*y{E�ϝi��A�*�Fh�E�dC�0�ۓ<���Mw����ý�0-Ug���i~x~ѯ��	����
;��""��FI-ѯv��'�L��>�f�ʠ�xn�=�'.��Yt5�9)���b��8��խ�n���,MJ�
v�P���㈳h���R�7ȡ���l1=���Q}WP&_2!2t���F�=-e�~�u�^^o�꾍��^ݓ���M.�3�R�:�r�ؠٗ�!�����Pم'�qQ������"��nwצK�e%�^�}u-���^������%�k�a�!�ˋ�|�}�{��:ؕ���������*L�h+�hQ����v��Q�;;��Q�z�ז�\�|��H�Q��\#�{fr�p�C��0�/���F��ԅ& C%�$<�,m( vd>����D }��>�[��s{�(�2���^��Q#q���{Ssŵ5�9�EmWЕr�WŦ+W=���R�t���k���I��cbq�)�0�x�_2��
���(�if�B�����'\2.r؉l�g�(�*���zߏ�Cm��M���߆�:E2�ѝ�m-!_I�!��M�H�K,��"�uY6���Ĵ8t�!�s����� ���E�rr���H������X\�1b	�<��n��8\1�\�_� �3`/[_����ǣ�c�v�U��d�l8ngv��� �y���n�y8b�i��b y�5��(b�N�\�RA���Z��`�a�����JQ�����Ԕ0�9!1��.���~��}�hz�ty١�TL`tT���I���*�e
)ҧz��Diy�ܿǉ�*���. �$!�0����fg�g~�-����d��3��g�h�Y��)$��i5Jy�?���Y	:W�W�����CԌdC�L��|O�������¶��_�y�⺪��}���[������lɳV���@�Ix-�*�oTD��yX�������ԱÛe�9���;;��Y�$C�J��9{�.���u4��8.����0��~�_����GQ�Q���v$iֹGD#ݥ �-�m�9vd��Zr�}�g���4�&�P���&�t��T�?��0�(*�����{�HB-�Uh�%3#�/��`����S]4�>�8c=5����m������f�h�(�������� ���ÿ��N���[L���~EI�?���UAۙ+�d��^1J�������y-/G\�/�I�@*�kP&�UF��ˬX?��D�!���v-�1�ϴ=���){6]�ڐ�"���J(:9fb.sHg�R��|���˸t-�>�+A�mV�.���[��f� �H'�`��m	�����w��!|�Z��:qT������&/&����,���Sӕ�5$"��z����%%���=J�`O]"��ѭ58TTi�K^׮��߳υЏ�A:;X��f�����*˜Z�t��1���M;KʊoH/1.;@\\KW���Z�X���c	g�6t�EX�ZV�&�*�D��Y����X���ԭ��<��S�Zn��Db/��P��U��<��K`���[BO�S�O��}E?o�&So���^A"^>1�֦�{�?Kc��3 �Xq�[е��7����8���Rel��`�BO,�_K�|�jQ�F�f`ɐ$eˏ�lA�4s�o;e��"�����a j-Xt���t�K������:k@�-��������rΎ�ց7���ƀH���ſ�����ut��+�RȷV~�M�h��y���R�U,�|at���B�n��L����R#�G}@��!��
U�B����T������Q�;��7wT��MJb�f�Z8hx:(�l�g�$�	�qfދ�)�	��1��#�Wτ��a�ccx1+_��ɀ"棞JR�RC|t�u����]�:�<H�h��u�A�D�i��j�m�D�A����^X�ǽ���yS픧]:Dlq�]Ov�	�s��<�:9ܖWGi��Y��p�2��C��l����6PU�Un�O�l�^\��ۀ.��d1�)��u;^��G��n��bϥ��|�����;������P2�D��v���хD#"�����t��r��?�!D��X((���	�Y�?�ŝeXMp�e��ޅ�bnm�8�H*�N�F����f�E+4Й;��f�^� �C�-��M�V��l ���|\@�Չ׷��;���1�n����⣈OW�(*ސ��@����O��@4�ucK�c�{����2&(���#�J�Iό�U�6�j�'-IjY�!�f�-�����A�`���v}�O#.$�Ď\�cӘ���@	*j�Bɪ��j�y*��6D|�"���d̖�#?�pt��Q	�h9�"L�PL�������~nWR�Gϑ_ˢ�	�	ۮ�P{���'nL��$�"�*�t&{j	�oqM��t�f�-���f�EN+V�߼���#��I��κ������S�yL��LB�e�����&�����*�����0��b��t�R�j�BWL =l��Rz�7��N�e��H�s1��k�z��{?�Fp@����JL��R��J�~�S'	�����-}�B5oo���~��_�{?Q��)�E���?o�8L����m�U��fs����EI�a�W�Y��Ч��x�%%MQ��}�.�U�P�W�Fh����(uǩ���ѻ�:��)��t$�Y1��Q���ԅ� ��3)�*�sg��2=���w�᝶)�!'�M�U=�
�HO8P��m��4%C�tvE�5��8��t���0��02|j�(�R�[� q}�Ӧ���Y 4�T���L،���QϦ���q&���6: ���G9�d����^㪌�jr�{�����a�z]W���6�+���dc}$��X�����48l�v�����Kt@�1ʨ�.t9vP_��~?��n���N.�`���y��I���6�ɴ���J�ŧ� Y[K��:={���Y��LP%_,�wШ�XbgM�)��h{��JXR��;p?�9ةS(�tY�vݻd��z5[z"�{�/��d���!��eshr�i=fb�����6.[�A�
�7y�*����ݧ�<e��d_��~���M�M��]D�c��)��,Q�ެ=:�
�H2+q�]B$�S��>��%J���t��tF����[.1C=]���!�wb��ci��Nr��H��im�|}�!�:	T�vC��}����"\���BC�;�x�ew�S�@3�&#����z.lw��X.�0�\+(���ZH˿p)2�`c���\�+�( _	C���CtN�j�3��s�u6��f}���Dמ����3��Ky:�6ٵґU�a�\@5\rD���q�x��}h�����>����KS��k6-o�3!0O�ʨ%��e`�jD�1n���k�I�9Z})�W'�`��$�j��=*�w�Lh���^����U�Zip�i�G�D�0�c�I��}bvm����<D�9c�f�j���h���z�H4[Aǳ��A�E�J<�I#��w<������C���D�����e���Ҩ����jT�R��5��^��V��k|�6��$�R_6������}3��w�B5��Y���OzS�.^gvdz���Cz�P둹13S�t΋��\@03>NYC��=�_*�]oa�%�������H �#�@g��?�6��6��c��q�;�}/��_+����ݱH����?_ �/��yF�AȆ��m�P��sT �� pI6L1P����,�MS�)=���1H��}ݶ0�b�BI�NǛ��pχ<q�׆��A��l��WU���D1L�F����Gp� �iW���o�
.��a^zI�W�ɀ��ρ-R��QyG��q�FϾ&4j�Qc�+O��	>�b�ckR��+��|�|���� v��m�e3��\�8
�Rݙ����Yx4�����sCzO�v��[c��@8`8�=Z�F1�yO�������F�T'fO��NlX�������n1��03�hL)3}����ם�M�f�3�WQ���잢"�����O8��-�M�Ւ�1�v�=�� �a=�����v�@�)
�����}�B��L�Sȋ��� �Rˮ9+��QxUk��=�E�� �	e��rߘP�.M�}~��fӭT�I5��rt�t���)���Q����9�v��JC��-�o�(����p��GJ�-<��B������]%+%=����h��K����n�"��;]U���5�l�73-n#��Or�b�_����q ����MKt@l�������B�"t�?92�RFYH��=]�/A�n�9���B�u�{�;���Uj�y�  Ë�ŨP�:���]���ATt|.օ�,B�>�
M�(a����q#��p˄��� Ww�,Uz%3�M:VKY�H�.G�G�~���u�%����n�&����5��6i�q�A���/�E��&�A~��V� ����_c qFb��HRj�O��#��ឹn�����6n����B�R�j�!�b��*]�b�z�S�DC�*0�B���O���{2�;�1�h���GMt��<*+G�k����dS#p��J�M���[��`?���y�|Q�2r�V	۪pv�`eЫ����'xO��pt�/�V����m���,;��﷤s�!5��&�����'��Y�����M �#��i$\Lt!�&�5F��Y@����y�����	��Kz��MBX�ɬ|K⠼��k�֞�XCP8�P�XT�%�rʾ�-��y�E�xc�5���ػ��#�gS�eb�/8�'���w3�aH�Hp-�|���T|��yWb���y�LD��1��ބ���7z���Y<���%o�γe��ab �d���a�$�FB]}��Q��8ԭ;�-�qy�i@e�o��E� �$�(�b:�0}Z�@�sa�Y_�uI�^�r@���֖+ݏJ���J�4��l�p��l8[08?Ut�)��Bi۵!7��rΔ��i�H���M(��.-��#��V騏�AXy?c�F�>'�Z���!���Z\l�������c�W���$@8���ɋ��S��?
g_����!dY�q%A�������˩cC��{t��k���VhEăh�@[5�@��ɟ�r4qV��;�����LOY+ i�'ҟsF��t��̜�`��8��b�=�K���a1��~�E��Qۤ�H�[򍯣��z?�:T�X�]�n�5}��%*	V۴�h=�W�&��k$�5Uj�|�����2��5p�M8�ɘ��@���C��Mf���
5��4mS,$�R�P�ˊ�8��Vw�/s���ָ�T��R�#F9v�|���Z��M�^µ��&�8KZ��ZN0*�N)?�'����'�J�8[]׵7Mr��1�L�{��1��~���:��� �P����c���'�ǃ�*iY�?����1:�}�ewv�G_iq��;���t��y�%{����i%x��Ȅ��� ��_��o�bv��u���qh^|�W4ӊ���b��	ӥE��-�ߡr&�x5�� ���@����Ti��ݴA����J4�s�;�G�H����tll0�5/z0��;��y?�=+��Txk�g�h���1�o���N�Z��o4�с&��-@,�V�U�\�Yة�������W�0ɤ�vu��q�NZaj���M�@�#���i|�4��Ԣ�X�>�~�J�U	2���%*�y�y�"(*�$�/x�	}�<��6� �Q����RT�d^Ǌ���&�w�&J�P"��wr*���Iv]Z�l��TU�1�t�F��&*���>y�;b&��/)m���<wa��}a�j��R?�	�{��������$i�٩�S�gܼ���+��Ú�jԵս�BĞYu{QW����,(+�5��l�S��V&P/��JbQ���yطD���*sՇ�=(xl�pF���|�%�tR�;9/IA6u�T����<��bQ�&5�	ua�h�i�Z!��9�l�i��C�[Vz��9n���I��lCGjv#�}�7��l���V���Ed�j5���h��=p/�-CsN�{����>Y3�U� d_&t0'�ƚ0@n��p���,D(�r��Mx׮�K��Fj�[˸���t7�
��.27?���{iKq�E���m����{Y\�=#�$�Z^�������d���ދQ\�FS�b?����=�y������5?�MO� .Ė�m�B�8-���� {����]�L���%�s١�U:�$;�g�d��]<}߾��HF�UI��M"~C5�ؘn#�Y.Pl5�f	��ɑ�x]�G!��0	�N�mVh8�#^�a:}H�9��no�z�t�*5���;�7��I��&�#�C��T�*h�ۏG!��"���d(�u�
�fr����g�B�@�c�\�.!�y������aL�j��项j�燚;�fM�i��'{�"HҒ��:#�'rU�j^ʸPd�R�Ʈ�mS�ts�N��K�t>���̌=H{Yr,oB[c�� �}��P܀�MjyF��)�ʘ�ELx�0Nx�j����lSIr�����ŃAu('f�զ�=z1l��&;5bj����3��k�i����Ѵ]���n`��TKC1�1/2]� ���Yv����}���ٟ;�6�"�l�B� �"!�N����e_�^c�Od�#�#|$�/��,1��,�����>�'����[��h�P�W<�k2��*����ݜ	H��AC�f{WJ���-�v�Ac��;�ًU�E����xө71`�a�L�tq[���#(a`Py&���/�k�d>��nL(�s���X��w��^��BXr=��/���v��X<T˃>�.�Z_���F�_���^���b�P-���	<�I�U��dؐ���t���0�r�GF�y1~Q�OQ){Ar��K�u�V�#r�7$��}�Q^9�]�#�R�8X\�������^
'5Z)��҂/)�^���r��;�hu����DD��l��i
A����<�n��@���X���&���>e'�:��r�gs)Im�J�g�~��ǓaL�I������՛b�b��P
E��}�)���!Yv!���w��׆�;�um�b���1[�"���W�4��%����N\�"[�Ӣ��mSS��i���OJ����"�瓜��Sx�߽i��T�o!�SUV�jWM:����h�Ҙ������%��Vj_�N�$�۾U����=�&,�%�9Qh�9���#w��:��'�OG�A=��A����KS%W@\�C�gL��� �1�ֿn�S_�w{j��$��� �@Y�Z�]��xW�&�y
 IF�d#��v�}��pٱ��Ҳ�L��l�*অ���hN�ѱ#�<w��s�0�Cj���|/�f���p�s#c�dx�f#88$�,Kl�bs��a��WWS!�m�9����P�"��`�d���GP����M�Z5D��+[�:�g>(�5��>P��qS���l�'"VҜګ3N���e�[x���v�S�e����d����.lF^�n�������p�x�i{��N���0l(�
���-ǳ.:���>�-����1p�:tȅ�Oh�UՇ�$�%(/?���?!�����3r��x��3��Q��xh�>�`Wd��lx�t���\8��䗎-(<�Gh���E9nt�m�n��U����b8�pbY��-XELu��`0F�k��� �D�q��@5�	-~����gX�� ��t�4�N���"yW��ܕ�5)b�+��:��8�ڙ�jgL�1�d�3�V��Jrye���X0���O��S)���j���@�NT��=)ʕN�ɂM
���4"0�~�5%/�kҕ���g:%`G�)��q	<kWc�W@U����Қ7>9��h�rHu^�7�4���h�`���?3���+v� �o;��W!��V�ӸHu����|R�pw�,�L ��#�^��k��4�q�IrV��QRW{���N�z���^Q�� T�?R�D�1��:�2m'��=��Gj�Wy��%$m��b���|��vjO?���������<���e<1$#Zo(�;@�'��lu%g�T۾[�����$%អ�n)ƻ�/yзíJ}c*}�֧t�U2��-�]���ۇG�����|VB��'�0����L;:�k�@��4���+�� �Ӹ�������0���hj�C�g]5u�`����{ş@��Hy,i]�3��F�2������� ׷n�-��[��c��S�	b��(~H��X���IVJ��M��ؑ2��-�Xi:��q�:��S�ȵ��[g��VFs�[��'Go��;��F�(��ܐ96��t�3ֱ��� �����8Z�}zP���(�
�@e`���S�8ό��%�-�m�����9��=�s7�{��bYcxYp��;�����Z7	����%T%�@�	�A,��5��d0A��p��M:x	����&b=Rh|ц\q��^a
(�o��}��i��z��}�P�l�5֛�x!+B>��~�7&B��0�~Dk-�
�/Fu	���gmwg��P������mx���`;�oI+�k�~�R
l���9����F9H�d���ڝb p�b	Y��g�UPMm]�����镳�94����w��^�Z���I~��]�&~1r����5o%�w�Ee�W�	�?3��y����%Ir񱎴\����5ˎ�����X�
&H���L�ր��O18K�\��%߅MI1Y⧬�~�v1��L�56��������i����l���U5�z��n2�J�e�P@0���Ͼ����O�a��;�Dů��3(ҧA�,���) �������48c���:4)hPtz���!�Nm�-%�y��>w�<ne� ��!����Q���Wm����� �����v����oC%�6��R����]=��">�@be�M�Ԕ���������� �p�싲E]K�ƠY���l�r����@���#�z�S GN�w�A��̸Ō\lt��jp%g�T�����v1~��	�&�.(6t�k cED���~�A���
�d`zh��+� ��`�Z�%�
�ؘ�S5ȑ�}澄�����m�.�(�ۑ4w��پvFɱ�=��BT� 4YcB����)L��)���b������p���L����4�Hb$���ՈBz������l�+I=�2�_;���a���|���t�f��8�J�)��=S�fo�%a!�Z�O������#��OK�@���y��E����$k8�nz*Z��wm/Ș�`9�� ߷�ym�6�ѫD����_��п+E|�^�ݔ(6��m��=*1��%w�|z��W@*���4��l)^g_��wX����x!�mn�է������0�(�u��t
O~��1��|�1���L*̐T�3�Y��Dޞ/t�j��L���u�X��B��oA6�[��?��ӭ׭���MO�^���@#{_$�3Y)፶�I�,q}F�pJ6���ax*�M����P\
���6�ɓ��?XRW�'�#�g_�r�	�����{ �G!Ԫ� i,�� 65!�[��mYx�ݫ�9��`�� !�O��� ���q�Ⱦ���%��j!�F��F�kwXu��}�4��6��pH��������VHVa�w�謽��jze�����`��*c�z�%�а�ej(���WR���h�V��P��X�g��F��j@g]��EX����Sѩ�y���p�h�O�]j�;��:}�Y
��~#A9{�U�@���e��>��E���t��P�'1U9b�9���1M�L/��Vtp���z��ԧ5��e���ѣB~�1j��-,C��8K����'�>Z�����М��b�a!�*=�y��<1#��1~3.r.w����h~_��epo��-X/�!G�9�[���aןV-�nQ�q�~���䡈���P�L��[νx��c1W��%Żl��DJ�['�2�Y�W�$#��b�m�'C����Vp߲m���E�e�*q n�rfr�)���V�3uDW;���b��jW'�;� �O!�AǦ�bdjo��y1�%|�6����Ԛ��
������$���=�h�����D������Y�
��x�^5n_%�"lڦ�T����w��W��K$�r�=�8⤁vhip�^��1��J���4tN
��:�`������:y��;φ�$�9Q��R����g���A�%���#��yn7���Į�d����3U�/2���q��.�B��3;T,
O�Iv1���MSb����k!.�q�ߏ��T�x����2D�g����x��6��]�%x��i�u�y,p?�	e�-�"�13�u?І�X�jy��:Y�,��ӴD3��6�N.�΀s� \;=j��Ƣ�l"�S�|%,���SE��Fz�O̺��EZ,���j�ΐ}�.g���i����0C+��Z!��t*v���8悁�ʾ�؈�D׽A����ֵ*-Nte��ήk3�vޏ;O��잗��R�V���C G-�=�\zy9�P�;�����-���XNp����rz�tǞ����%8~��KW�c�x�D��2hܝP" �\�/M�m�1��r��IEnJ�&��#�P�w�����a�N�������C�Kȩ	��� ��NZ;�74���HĻD������yL�^�5)�Ӵ�V�K�P���=	#ԟ�0rB���r(\��sc��/�5̇��K�nE�7׭|��x��>��e(o��e�����z����'�&��)�bd�����Z��0R$�"'T�+�����W"B�`b�k�l�/\���դ`� �3�N:�G~N�'����{+�$���1k��Ǥ˯��Է�{�LZ�4���\����Nbpu���V�Ρb��#� ��h��s�f/*-rp��h\��������v���t����O���'/Jt�9�O��ڼRX���KK���j���h�Xw$[���:�[���w)�zk@�p��f[��:܄	6�I�����0G�9���xi�_�]B����9@�̚p� �aaѺ�\ؾ>h���M�^�Z1@����(/�Y��SR��(�f�=���TR�%�h�������0��Yȃ�T�f��ΡĞ���a��X��)z��-!z��8ls�Ŭ��yXm�՛?�w��u���(Oz�:�����\.Be�`�T�y�v=}���&9�G���q�0o�����8�bn�r�C,	8��ֹ �����/u�|�f�y���R������J]^��s�D���fN�L&Ƽb(�{zKi(~�>��CѸ2�[�5���P�-���"��9��Ξ���#����g��fՈ]!����[�u|��>���I�=��A�ϥ���6���͋[��N/ͫevS�0B�o]�|2�;�B*-T�s��
`����|��?����p ��� ����be�eBq�7EJ:�I����3L���~B��U�TR��ے*m��@��HA���yQ=BG�o�8��Dߴ���$0�j��L�}��)�m���%'Kx��y��}�)w�n<�l�O3��<�q.i^����� n����}n/n�<y�MQbb�A��0IbOC.'����i���Ǻv��<Hk�����Ut3��'�@3ܑ��ꍀ)m3}^��b��_e�s�܍<O>�w�?.v��p�h��Bǋ!�mHUE��k�>_m���وt'��Ld?�:���1-�\h��W8칣�jG�Kk�9I��E5�z�����w��>���d#G��Dk�ƤhB5���+O Q�qث����"c{['����"00�I� ьi
�,a�p��;�+��b��7�{'�QR�c�Mԟ�jY䄕���U�fCQ|	��1W�#alVHWA"U���vʻ��I��a��,��� � �0"��R�Ȁ#��qǤ���<0y�֘E����- Rڏ��唾�5�2���r �Qb��~�+��{���q[Uxп'���d����2pQ�����ժH�k@�V�#s%Y/�- �y��N/{��[�ZW�BG���yw��1�}�'l
������A3{�L��`��1��u�ʸVg�/J:�b���|�E��ŗ��m�!����(G6�и&�C�X����zz�`��w� ���'I�a�SE�Lԉ��7�-��1�в�H	�I��ߧ��g�y�|>;?6��<�B�+h��8ٍ؁��Ƀ߲�����0�u˻��y��*|��d�����z�A9�D^�Y���rÃ�?M4I]C��m�/v2�m@$p��T����D���̔��E�2ro��1��N�9�N�L�_�d�|�1�W0[�u��0�rRQ/�H���"����%�� ���0��Ѽ"H���,�	8*������ޅ��};���i���_�����B����P�Ŗ�J��<���@sZ�$����xC���!K�F#I���)JD�RoKr0��! ބ��{8�f��0B�ț��6��Q���#�Wy�O��{��J��>&�������:^P�|s��s��_	ᣓ��&ʟohW�����fj���E�?#-&�b���
��OIO!���;]ULy�>F7�se�D��Wp��S�k�P���%�����u:��Y�F�:&a�D!k�n�&�(pEZc`��aG��vn�<����)��5<��DJ���N|��,��B7�z����
���Q�w��� ����f�B��uK������<����@zW������z����]`�v̺�c�XSUr���86-�#	-�yC	�!'�q
�PyT��� �N�w4&��tmx��h̇��Q�A�H�H2���:���ж�e�Ö��}Wx�����j
�d[�D�t?n��	�a�=��EL�g�!0�f�-�����8l.p�l�oP 	����']վ��I��ւ"c$OuN�s������_�B��++&r�E.�v��X_��mAO�?�>�nK���Hj�={	��^��g�(D�=}Q��(+��p��Y����C5�9_E8 �g�,#puT��of^hG�Ǧ�>p��5܋��.�*�w�k�ݸ��5��\/YW�/�ma\�n�8�������֐ϣ�݄�!�d�O�i{�X*nnĜ�=��I�� �����iο���n�����X�� 2DV�4;�P�|3K�����5SW�5
@�K�R"��ܘ��B��"z���J�Z%qڏ|hN]�8q��1`(I�<d��@&J���2�(ebޕ����}�n�M���1+�]"��lԺ���p9>]�����2��(nP��?:�f^��媜��ɜ�R���щK`^!&��̑w�BZ�^�g�!��𨾿��)�[��� uѿ6_ِtu���"��O��!�券���_�n�vQ�w�պub+�BL���XlC�G~�n���P���ؖF�6�G�~$l��t�7�wK��V��E?s���h�A�>=�w��"�SGRP3a>���
z	�;g~o6+����I59�����v��8���&g��s�%�G[����Wα�V�d3ZX�T�XR9�;�3�^eVE�m1�kGphfL���[ԫ$
h�F(�D�R���Y*�Sz �t�lM��%K!�yL�b)�دj�-�-����E��$���_��9L�j��D�t��6��_]�(e0��"#Uշvɨk��Ǿ����tC*a�7~�.&���!C����9����oFpm��w&��E� ���.�	q���&`��b��2u��U�:G6:9��V`�*���y#�M�O]Z��G�r��W�u�B��O!V}���"��/�s�0L�I�Cߡ����|�����MH�*4	FO������?�Uq�6�*+j}�2ȧu�Q�I�,�''��K�3�W�oh5�@*3:R7�V���MH�kA�3�ˍqt�&�5���w�)z�J<�ڦ�+\�G8�3�˯�M�s҈2�$M���@l��t$Shjv���b��<;�%�-ٸ�)?M�Ʀ^Q��nA��RS�C5�TmCf�k�w��:��ģ��iQ+�w�3ŷw�Э��#D�F�H�[H\�D	h����/���-A3p�ѷ�Ψ�a^��l�FO��8�%�c��F�0`u=:�/}qbW��br-,����O�u)f��:F��^�cz1�YU�Kv��TR�d]�[���'MT0y-G���� 	uF���Ɇ��R�ؼ�m��0�ҏLzɱ�|�����z�g��PW�%���w�ر-�:VM��oYE�_ȭ��VE���d5a��˵/Z)[���Pč/77��rC���U�]o�F��ٜH�����d�۰�Fd0��0ӓ��d��b���*_&d&)1���hQo��e@�ۻ�sI�0!9L|��.o���N�u/��n'D�(��/hm��P��4̬ɽn��u�mT�A>����v9}�b��
�d��7ؑWz�Vz2��2qv��g0�xO�"��3��o����#
镉l���3��u����`���ٯ}�<݁�I"ԍ< �(�Vw֜5y�gS|ݿN/-�H��N�4�GBS+�aMW��l�)K觮��8t��vU�v�)���GE+�O���s�E�Ar�5�uuA�U�|����ԫ-Zs莋����T�`p��#_;��'�ˊhܱ�6k2�&&ҠHn������nյ*I��L����QZ�s�K��ㆾƢ�s���7����e"nc��z�����{��3H�UR@�r��z���.��42�Q3M�K���R?U��U�ݬ����U�B���Ԋ��5��;s���	��~���ٲ�JC�^s��� \�G_�3��^�[?�:���
�����}BU�v��v����cz0�,��32-��-$�b�S�_�E�S۟����,��j8�k��������ݫ�.�F��m�S=�5#��ˉ���� d���η���]m����^C��a�u{�@+��n�w�©�H��"h�dɊKA�������>�OҶ����/�B�,����1�X�2�X��R��:Y��R5�i�r��#�N��G�������dc�
��l+c���~ڷ��;�\# O��p�i��z�3�}���0���K����٭��1�(f�߮s���{�����I	�|Bf\ Q���Y�
D��(����t�K���l	�݌��{ �,�F�
�y���>���	|���gE-�}"%�wm�x�����y�G8�D�G5��R��9�՞���BXs=��ԭ�L��+P��6�.y�p'`3�/�*p��B�	�X�b䙩�:6�O���ă*M�Hr���"�`�(����d�/���dP���0<%�ꖁ�x��֜o<de�2)B?���/����n�վ.�	�z�Y;�[��V�m�"�I����2>��(�J-�������%��ȼz b�lJ50�K��2��8�L�f	�E��̶�3#�� 2`���?P��҄w� ����'�!mc9�;"���2ȟ���h"�ו��U'�T��R�+�h�r,��$l�ﵔV�#������5,g��V8��yJ��$&�]��P��y�5G�~�xQ����A�t,nAZ�gU�Bh��D]����7y $��}�o�S�������%�^�g-�ϗ~9:�z������ښ��슷�2�*f�R���i�ÖLOf]���r����,Eᩀޫ�>��+D�"��iyְJ��h�m]>2�Q3��%w��?ED8��,|��������۾*�CF`�]D�h��`�dv��υ0@�6{��m4	�A�%��$!).2���ȟQM�g������Z��ᾴ�8������Y��5�|�y�:P�5LF�'*��B �t3�5���c 5�YZ(������cbA�+��D:upV>�����:�=���u#�S���ߊ�$�7�o����ɥ|ՒMT4.�gsm\Z ����,#��D�+FE&��G A��=���謶-O`��P/�im�ܦur9�����c�X́�_jj��S��Ӯr7�=\�	P���7��ݩ7�\��o(���v�/�@�_a��w�e��2�HT���-#�-bZd�s���`�X`Z����9zis������p�Ւ6M6��n�Z��޾�������L�%ߔؔ���Ac�ۿ���X�[��}X��W�e�8�P
4�|�,�D[����wE�F{9dA���>�*6nh)���͸粥n�$�tc�p�r�VAM([֙zo���/�*J
{ezuP	`Q�j�		��G���di5I���[���vd��n�O�_��-8iynq͜F74�XGfr?�!L��moA��w���]N����7��Ob�y�k'ʷ�������Y�?�����ڢ��g�$����lWo[a� ���:�/RV��ᧂ�ZEM��ח-��45:/�C�"h\̀y�C3��]\�Ɂ�v��N_Z?ȃАs2}7y�_�t8�a��O]F�8�MM�������[���#Ztd��Beۧ�f�!:����]����1d;�ӯ��/�)+z �+h�ŎX�7�2W�
Z�d5�Qs�4�����}�2˳��r�/�l�x��̋�F^�U/�3hB>y�~��,S���P�Hf�;�8k#�>�j���5%Z��4>�AC�ff�}�X�yug�4���3`dUy�|-���X�ZG
���v����7b�)�@ٛ�+cu}��Yr�!-J?�$ܮ!Y��h16��]<WGX?q�(��_�h6l�l�	���=N,�c�aʩ	�f�=�k4H���3��.�xa`���7ϑ�ٟ�#�2�(�z��X�.��d{�u�<f�t��V	�Z�KZ�?�U+Џ�+��'�����{�/�7���c'8���Hx���v��V��|��4����8�5 G�C�}a�,ڍwtMhUc1���6��p���`IG���'ۛ����<kV������������|sb"�Bp��Z�ܬ26�tƉ*ž�s\;(E!��]T���_&~ȹ�{l5h����^���YgФ����L-�ѭȹ�P��"�{)�`"O�lm�D��l�'6&�.���0���:L!�2Q?K�\���9y-��1�{"��^�(ᨠME��_�?�> ��ͅl��@w%&�23�Dʧ!�b��y�`Z��Cd!b/d%Ʀ����T��m�V�^��T��}�K��*1dR�r?v�1A��n񉦀����~�J�{W�#�o�z*��C�����ѓ�E#P��6�)��M��Z�_5m̐%�aGio��Ɩ�o<�O|��(�r+*QP��_����a�{�m�#���Kg�7�P��c�2O�XZ���J�!j�;H��=�����w����!P=`���+1����Ń���i�t�48��� ���U�~���#��,�AJ��zՙ�� R��e E�zϻ�9�lW����P�"�
�	;���5��wt=�m)I��߱�f��ݞe��*p����A
U"8�Rx����o����)܉���<g��]�\38�08dK��]0����X������ꑐ����-�g�<�C�|x��$���s^�_Ǖ��r�y����kѪ9$�$X,%�D�`5yp��1U��"
�^�Z�E��tDk��Q���W&�)L�0!d��ו֤o�2I��I_���Q⛞�eۄ}���a�jq�K� C�x������$��O�`ԧ6�?���B�;k[$�	���O`�~FN�$�hmѡ�jU��ƾ{럨H��km� ����5�E��px���S8�{/>�M��E�L����1چ��N4��u���Y�'�uY�/v�~�v��W��5�2b'��,U�������t���U��d���n.!1nMbvtl<2� 9��L~8������(JH�S&[����k�4��!	��Bψ�v9���j���D�V��#ԨL�p4A,�������v�k#��l���^W�7>>�>}&m{���ڿ�$��,����^l6mթ��y����Tʯ(t( X�:�T�V�2"��7��/4�#h���]��F�`78���O ��ۄ����&(�	Y����Q�N���^��J�^���K�Kcܖ�R��wI�p~-�<�64�85��O#"�BQ��T?�y:C��(�^���s�82t Z���z2J�t*6[���.�=<����mK��Lɞ ��m�K�ib���?�I6���M�����W�G$�d���\�g��|�G��r�|Ñ���L������͸�r�*���=^�L[lf��-�s���H��WΚ��k�u�룩S���K�
��Wʑ�@`��"���t�@Q%W��+р;����md�ؖ�"lp#W�B�����U6����+D�b�K���s��%�7��ӗ!�g�S�S�݈���ϧ>�"a��%�8��}����ڤ�G���d�7�|y�dͳ*�����ci��/�U��)�)Ԥj���n�A�#�{��hՈ��ۋb�\�O���ɬ��ϰ�5���?6�[�l����_�\�����&�np��3�������:kXl�E,�Ъ��5Q)p�ORt�O"��4Q����� x���Kk�8U�qVjW�P�:Z�)���u��f�)O-]����f*�yj黰�RC����9�!���mW!�(��4A��0�r�������Z㍩�=n
j�kc�F��y�C�\�e�*2�J�+���R��p�xc��s������(�3��K%�:����*aW�e�(�D�Ԩl��-wI��|/��bm�>|��E�u�̡s�fո� cՕƨ�FU�_7�~���fw6�H���Ga�t�c�qU[o��V��Go�v� ������o[��R�
]�Z�t�M�hC��eNI��F~TvL��8i�!����l�}B�����O�1O��Q��Mc��X�@��<���!2�h�Gi���H���D�S"�( �{��&�Z���}�JS��������<(�|c825̮���9�<�{� |K����\J�"2�/���gpFT.��g>�ib��ج�ufu53.U�Ҧ-�A��[ �L��ȃ�UY���xo�2��;v3�b�TG슊[ ���w\o�d��r�);�֦�	A6­�vBՑsb�6�V�%\��	Z�m�Bp)|�&F��b��,��h-+j�2�k>����
@��˪*�ڬċ8}��+��}�����#�H��PWG<n�Q�T�PfC%�,�@��{�0Z�
�Ay�p,�B�
�FzC�Ðra�DH-�EKC�oȖ��h�IҾd�fw�N��<q�a�t)��ci}�INu����~]�UW*�C��0�Мm��{E8��IRo�Jc�V����|�	R�j�n�}���7dH�����Z.���i�N�@e�L/.O�3)�����͚Ř|l��}7xXC�Ӕ�����>7�礣�\\)4��|�����D�q5�r�l�ׅwi�gƚ��soC'�����6�-�ܲ�1+��9k�Pw6[n�[������w�&�tS�0�I>w�Q>�����(�~an�ђa�5��ʄ�5U]ὠ�J����N����Gv�R���C�׋\a5�t&����s	�-W�_�dv�;�g�;4NVc��	��	�5;��̾���%�	I*�=z���P��6�M�P8j�'�)K+�gM��B�LY�?�װY2������
%Ƹ'��,�>��_2(<�IF��n䚫T����;/:N��i�&2uǿ1I:;��A��Fn��>��8#�� =�*�7A�:�.<j;¯C�,�Ҳ�ũ�z�-ϟ��h�C\4$k��re�����MD��z�U��A7?U�P�K�m����SK��n��Q>���O�`qVu�ʬ4A����3���$��G�$���6l��%�X��Oq�_	���{�V��w�ϙw�#�+��%�-j�s��!��S�!$�>:,;*�N�l�K2R�❇^�\��"Q���7��g,
Kد��p�	�*�E�ܳ z*K]��ji��ɤ��<A�5�X��d��ep�Yj�H���ָ��v��Yy�^)��R�|�1e�
J��怢�1W/L��Or�����|��)�9��<���7<HrYK�&��Cw?o�F[�����=�-mH*�l/�A�%��oT����e���,�������o���M.�0����Z�g�[-���e[������ݹ������s��d��o/�h;}��Qo��
�O�ԕo����>�@0�{Ź �s������R3@�:����7{�b��\�2ׅƿ��cm�KGRK2�>t%^n=�k�� �Ab���,_Փ����t7rE�D�QQ]�9(��{�Uay��6#ZL_�7�H%����~��4�V� B
��#�Hc ����|����a�ia6��nef��n�uS)�s�]���5�˥κ���v�:'z 	k��{����&P���u����[����Blߥr-�����X$y&�������B^�?���hHr#p�{!���L�1��	�̀C��Qo&k����[P8��z*��D���K�7{���8װ��y��������!���7��"�cz�5s�o>:S���f^Ͱ�5[&�S���u��vP�8�[T���a��u0j�%>�*f(���	��+P�v��kR�!˛8q���D�^]�ӁI��>�W_�ï#q���Tk_:��|K)�U�Kь���x�M��Rs���,����QZ��B�m���,�`G̨��v�:���~����w���`#�4`6�3� &���6>*��f�ŝ�1��![P5���d^g R�8�iYj)V���X���Q�����2���ш�N��4P�qЮc%^l8�t|��;��k�M[��4�z>�*���R����?�R�f�u>�@N��
�Q��#���.��r�.������2[��i�fx��2�vv/�����=<����<C_�ޯ��5��]_��׌8'K6	9Ҧ��d^��,=�� f�O7�n0���Iÿc�F",p��1��.��SIxI]qwno�7���X�a������u������ī��+��w`�:D���)�e;��b��N�+�e;k`˶��>^�7��
sgo��u[!�;���֏\��- �atU����Ef�0v:Z�����ɲ�ǻ�&pL�S�(`�#�T@��j ŧ}KC���{`2>�1 07�ir��Q�'gK;T�ܽ} �DL^z�hc6"���Fx|�������-]��d�ae<X�ZPX{�l�ѹ�;�ߠȝ;L]߅���?��o�\gV�<���I%��ל0��'�'ϋ���N���e�� Pt�J��p^LZ�|y�Ʊ��MD�8PB�\�(��E��h!��F:ǅ�[�9����N�Z�(�ʌ����'���d�T������L�Vс]����3>s��2X��=_����Sc��2�A�nLXaD���s�7i+���?]oس�Nb�Tv�S�GHk�����-�1���d_]hn/�h� I�E���3I0s��V��n*4�w"�BĄAQm_J��xd:�S���ץ��鵳cC�6װ`��U�V!�ms�H�šq�bv"�i2DH[.,�i��DQ�M���u�{bc������e˯i����J�� &�M`��}�~ ��5��aF%�v��� DZ�-�Iϛ�}ΰ��=�Fvt��y��w��#�u,��M��n�����ް�p��&t�;;��$�+�|��
�IX���d�+�=�s*?�+�#S�޺�`���	pO����z�R�4Ol�h|�=>�%.�yr�d3�*ۼSz��"\ 	*p��*�����W��O'�Rv9������iѕJ��#�'2���:H��I�Z�5$���>�1>T��	ZB~�"\��}�{2<�^M��	��/��q\L�fQ���#\���6R\��EJ�1�N@sr;=���#��n]D�8G^ �v�6�R�@5m�,�lG�>�"uER:	�[6���9�i��0/�v@>8���}es�S�Q�W��&ʜ��LnEޕe.��J����m]��#<"jr]�X�c\�^���6�.�����;Z�*j���y����>:�=��:p��,]�� \�T���Ē������B	P�Ĵ#`�r��E2�2���$y7�In�V̀���01�cc@~���T;ʆ}��B{�1LҍoX-午�]����hDߓjU���l���1e�I����\lu��fnz�J���~��4�׵=�Uz*qY�_���̴�_��K��;b ����I���L!�fRiL�|���fٜ�2WXId[c!��!|��/��4����"�Ya��hR��<�Y٤ęȓ =�>[q��s�6�ħ:N9�ix�����UbHB1T�$����m����T���FַkԀ5�^D����D�5@��r�.��آ$]*! ���r,#E�r[��XɊ��/�kc ��E���������Y�pr�&�3�С�}������)F���)�N��4"�(��˯з��g, )�M�y����T-�J�o�	�����y뇿�
���^Z4q��T}�F�);��~�����4�d�����%'�@ ��1�rE�{�X:a)ŀ����V�k;����`��4�]�'���D��KM�nP��?��L9�؀���k�q���˕����3}
g"������,t�pUM6Ё����?�o�����.�<�q�Nz�I@�g>��≢�]~[��0��*�U1BĞ����J��<�#aH��M5l�\�SR�g��m2N;��� �1)�5aD���%�?��:�[���	��A�;]����:k��4ˈ�7Q��V � ����1�������O۴N�H!�k�ㆋ6"�=����M����F-C��J��;�ǌ���1�<�[�$Q0���<�	z�����J��rڶ��+��ڸ�g�7�+Gf��:E0=/~�'�+���z��E�����Q�t�_������#/��m�/�����}���̾Eo��õ��p�������0:�q6�3=�~ӣQ��ap^�ﶨ�\���	���`߼�	�X'Ѣ��(٘��#S�U��O�����Ц�|`�E�A���@��ZZ��'�p�KӲ79ƍ!�܄�9J�L�������Vg��@���*��������s.!w߱܈��f�UZ嶲�����|,9����
�Z��"`T��c�������]��>�F��[_w���u\���.WHא��+K���c ���܌<�b�}0�S��/���_3 �6��"S@�ݩ�����;o��LTN�
��J�ְwh����}�PY�Ͷ�^��d��m�
!�o騬�!h�-����H�>ԑ�U�=��]�(�h�U� �aB����靽�A�O�"���B�6_����ʵŬm���Oy�u�X�̎�.3�ӡJ:�怡�`+���uHpR
9�M>'�l;��^��]qSV"f�(?3�m��I���+6@-��l���Ǿ��� �VY$� �k#�?y9Oc��P=��+��{c�@�Ŷ����z���9�tj8;o��w4Lԓ<�����|i�=yM�.C]H!�u ����9�u�������F�A����	���ю,�m�٠.Ӡ���n���l���2�no���������Q�9���7u��Ar*�{[�- �Ug�x���kĔ;�շU�c�A��_�La!�GM�����f��Q[�.xw~Nr����h�U�7���W���\p+K���fd!��Fn[�~��R]v�G���;�s�	�E=ǒK�V�K���YX��7�Y"���k�w��Y�я�� �񽈶�rt;�
/x�V�M��vx�uL�oCo�|n�KSע�"��u��K�8g��L.� ��X��e<�:�r���7zy\!�<�y�*��&@^����lZi�<I�*~8����p��$@��\Fd��;4=z%��s�2�O+\��3(8.�.4h��X�WU*����k��X�e�a!�p���F���p�Ȫ��`��������A}3�Lͯ(���<H��Z	E�j�7L���!�HbY�%[+�aʔ��`�)��i��6�T�צ�W���{L�G�o��Ҩ��k���j�v�����rx�w��.1(=̺
������@�pGkoِ�{�*��q#c{��9��T����J
�;;�	$����7�\N-�G��.��;�*�,Y�O�N�#`��b�P�gE1a5f�~��TǱ�SB���*� ��g'��A�	BD�c�6��O�%�ʅ��^-���y�h�������E���v�ܦ&�Z�z¶�dj(��	\1���3��ǲ�>;"���,�eR4�P���r����*b�(���;@���Mia	��X���ަ�&����$�4E���h���XD�G+Ğ2�E��N�)%?Qg)�� �|�v����*�;��ϫl!!�--=����q��ۅCv�ހz�h���!b?����}��M�X�����ur��MpgM���Ǟ:�}�/�8�#�b[�G*���+\R���+ޚ~�$瞧�j�p�@�0���=iJ�xߍ�;[��w�a'8_Ch�x��P����u0g����a`yNͿ�W�Yi�3#������pS |N�V"K�~K�/�zu�O��n�=�W��D��찹�[dY�-�p�9���>"t�~���~���)$q����+�e��+QW*�2U�����|���Jd;��:<Tm���ԅ���&�پ~��&A4�d�(V����뛀M�^��)p�V�O��4(���h\���-�!������c\ݘ*����)jP2�%� WM�fүj�+��Bvx�r�$�EJ�3���G)�8˪��6
�D$c�1���j?�<l�g���z����� ��!����d�Ii�\�hfy��<�T�χ�dS>�_�\�>kpUreBT�r�ἕ�F`�h�׀�d�A+��ϛ�������!|����Xπ΃H��5b����o��<g���MJ�&���od���y|�r��?�(��ӹ������v���,��UAC��L�0\�e�w�����$:���rO��ӈ�aL�\AZ|O���xۣ����C��ː�n�
�hQ����K{XO0}{��^�r��BP� �Й����m�hz��.A�������|sǃ�y�����{�?~nL�U�r��	QJjj�����U�/���;�y�l��n�� ��
8/�|���U�{%t��p�b�N�`�A�����bx_��3�n�c�͹Ԗ3��:�faA�	"�Jr�㼟2~sJR��(�r��ښR?8�Y�*_e1V�b���?,ه\�� ����7���~��Dw+X��6�|8Ǎ��g&^U[�m�������l�2�9��4'�Ѱ�þ&,aH��")��W��8���,m�5�%M��y���&����
�� ��M�F�KN�w.T�	����.P��xA�_�?Sg�4p���2�##�z����@�D �Y��`�L��X>l�-'X0�!^mx�o���)��(�Ks#]�"z���Lγ��#}v)Rq��5�8{빽<�$���`���G�;FM��#<��E���%ʊq��F��:����'x7d����_d9�D�hJ�t� ��͆�ξ��������WT���@!�bT�(ʱ�Ep��y�Sմ�c��j��th��l�M~����I绬j�C'�aѹ�d}����v� �����71��,�$9��.�H5x@ܓ	Q��U�Ӯ2)�jJ��IĄs���Q����B����irs8�� "�$��$xLΓ�,���atu%���m�P��J�2I�I,��s�t)[�:ߜ�Ε���V"��� e�h��T��Ju"�I,��(��N�>ni��K�\-�u!tȦ �.�#��R�rBmf��#cI�@���Ȳ�9:��8��Ȧ��­��Ċ���-8����_v�S4[q!�R2���#��Y۫�;{��2�E��~���.���Q�e^�+9�����C(<��	=�=�22�?֥FhN. vr����z�б(ڰ%��%+c^N�ra�am��V��g���W�#]c!$Ĉ)���p��# W��^�Z���F8Ik���t��ht�p�u������7!0��olJ��Db�;�潨Q6߻�-9�p�n�<�Ƙf�R�+u��C}��U5�3Hɢ�В�B����x�,����G� &�*���þ�h�E���FXA����ޯ,xW�>4�0�����gE{�X2�`T�<���U�j#�-�z��h�(���еO�����	��Ƿ�7�j���d��c��>��YRFN�c3�d�|m���vYV�.Gl���h�OKO�a�S�9iuf��U4����V��3���j2��Y
�2'sme�A_;4K�k��KD^���#�^pdU>Av(���Q��ac�y�a޺�]`�Yy�$d9;Qz-P�}�QEQ�%6eo�;<��c�2*�\/�۲@�M&�v��#+1�t!���'���U���W=�%s��2zl���]�h��9+�.���o���.����I�w&�|���]V�\n�m	I�� ��iӴɿ������3f�r��y�B��w\H}
�"B���yA�҉{��6 D����"(�����/��YFʊy2`��^�w���)Yz8-&u��5,�Mt
i;�i%�^�r����=;��k�E�i �����Pβ��p��>M=�U+Y�I�@a�שׂ���ß�bO�3b����2e��&jnsf��1��繉��]W +Gy�_e�3��'7�������L`A|�c�} ���`,+�|X/�O94q�iP`���x���|L�^����:��)�8��+�a��/J���7NAy	2�!�4��8YM�K�q$�j$8}&u�?b��0���_y�~��\�8�F=�8�\�V�Pnw^�Г���0[U%������A�����Hnk�uѹ�8��/�� X�oy��ZҬ,K2>8x=�w�)���uK'�ׄx� 0�ڵvs�_\�ͥ�	$svd>�	�d��f�����MFZ�q�9-�7�F�Q;l�'�GP���(%H�!�ǁ
B᥂��� Ȧ�
�i@|�<!r������4i���f�j�L�Ԍ�]��k��.��:ڤ�y;-4���A.�"����`���84�l��Eo�p
$��?ǬU/>����M����BN>�3KG[ZP��#6�R�ux`2_�d�ϓ��)��&G�Q"ʄ m��A��Ƹ���R�h��P�\�"����ps��]���U��M%!kR�#�yХ�LR��'[�kv{]w�����o�]Ϫr��@����'���`sy�N4�]�1>��M��뉬�<�'כ_���t�W��3cGQ��˹�-

��Q!�ޣ��Gܵ�B���[�Z�����%x�Fy|���F �<7_�ַ7��v��sy֗�n`��^��}&%#Ϙi�����4g��`}�)_f<��A�k�&p������ٱ�Q�YT|��a'�i���t�����H3�/�+����PV�F�36�Oyj��*�ݮZ�y5ė�T�/� <1K���W�wp�(jhPA3�~��Et� ��-P��3	��[�k��U�����l(͊c�Ƞzk ?��m��M����8���h.ħ�s���z|[�W�7A��ҙD�\��~�M�tԘ�ʔ$�$� n�5�͓��T���a��ު2�ƟV�~9ΣyN��TB��4v��i��i2�(�U���oT����;��zڧE�o�<�LS���40K������n` �6��j�/����k�컩ny��=oݒԷ*Dw�*�׺��~vp���`|[�I(�^�-������A֕O3s!�7�.�U��\4�+���B���CxKx/i�++3�'M#R�Ac��G�����)��+ßD���FT7��~\����\%�~�k}�p�BL�Yh91�?3��P�S�¨5Lu�z��q��)�Mi�<�XP2F.��h�f�7��Ao�]:�;��I^�!O����A���*�,�f�7Xo#�P7Z%)�w�
��@a�5?P�rCks�o��o��1(|-�+X�q�=��I%���2�-��|�[��kĽ�Zg"zThr���A�=�e%�,Sr�3��,b?�e��@J��y%�,e�e����C_+1wdR�Nf�~+�H%�C�O�(���N����aפL�[��TN��%`�dU��/�Ѵ� �@�v�--߰f�?�ϱmW��sa���d9��BN�Ә��Ae��X�J��ʢB� v�__��|'@p0�D��,5X^���5wJ�<oR߫�n9Ez����<�.�L���Zu�#�'|��b��w��BKj%>���1�U��}mf7�)*37h�ȍP%�MD��U'�(rG�ʸ�36�	mf޴n	����7��Nm���Ǉ)����f ���|g���1҄��U�Z��8fKz�L�}�� ;� W�8�ef$Sӆ`�)�1�3�!ٮaz��m*�����`�S�L9�--S1�NU��
���e��E�sp��#~x��E��b�J�jw���������]�a
5M�=/7�|�lK�ؙ��s�X�!�x�B��a�òZ���C��9�����n�j�-��z`Wiz|o-R�oX�c��ӻo�3{�	� ��SȿU���|�[`��zt�!`QŰ\ŝ��Bk�u�v��j�G�;쥕 Գ��[1���ѱ}��-ֹP��o�\tsҿf4a��6ug���\z�s��t���x�z��Y���ej�@�-c��ͭ�"�	ͬ+T����,�ޟ(Sd��L��=!�jڞ,o�MFf���D7��,�(��-��yD�ȴ'��v|��Jj,���<V�ʇ( �I&��j��m�u��n~*�<T�9 �Nw+����y���|��a�'e2ҳTK�`�Ģa�-k�o��g�O���Vv�Y��:q�q��� 1E!�c��dzq<�3M+�Es����
e��c7)�Q�;�iSG	�F�?joY,�r�M����u	�(�Jr�1����l�{�&*WQiۑ
��]��O�� ����[��>����b��{�Y��T�ˠ��AC��w F_�䎌����h�_M��*,���<�>Ҧ(pEKT?w�k���K�ɰ8�b�M�j�Bm�����s�%�N��_=戄��2��0�{���rc��'"e�{���¼)W��dR����?t�V{��������p*/��>"+ĉ3K!|�36���)pQk�G���!{6�r:Z)	L1�;>� �$0�w�5��~M��������7�>{��\=�h�!`�Z��]����ʌ��j��	��jh�c�I��}�1դ̣hO��kF���_8�]�ݱ�d��ZHj04o�ᑪ�8�d��t|����i,5��["ݓs�@�*�{*w�ZW���J�-�#�[���#t�،�\g=�)ޙ�T��n��v(��w�i���_��rL�kv~�qo�� �(*1Gbť �	ẃy����z���]���$��� ��|;�S�I�46ZFBȵ3��浕{e+���M��R���r*L$� �z���)�6�Y	�Ԝ��G�|����ڒ:�V�iu��O1�������ixy!��G<��Q+o�vL�ǅr���2P��_%��k���9�V~�i#:���ƻ�_�;!ETg�/���{�r��^�۲j)�|���\yr[$�����}jxnb�ŉY�vQ	{����������RI�*���&���;��F�C3��Q��� ����ʚE[���+)K�eI��0Ф ]���!w-�)�[þ�=B�~�����e�a�a��NpE�Q���=���B{��0����o�޲�B�*�5~w5����ӛ�
}d�T`!�er��#�`��!�,0���A��ler��!�5�q�Q�٪r��t?p븉Op��^?�� J���+��#7�{��i�4Yl������1ٯ��pܼ,/U*�xl���K��C���mmWz��� �f��%kМ��M�"��P�h�:v똏��-������C_a���o��z~'�\��V`k8��\
��e�p���� |�����/8 ��P���d?8P[�R�a��O��Ax^�� ��X�j��;�����C���@��������˫)��ԏ׿pz���Mq�n#��g��q6�Yd9;��E���	�q��
4��1=��[�����f��wC�%�q���t���GՎ��DHPg��������l8,E�s��"���+��~b�3�[�w�t�m��#��Y�88Wk�Oȑ� �Y��5J��SM�	�В]��I�Z�#&q�չ��f���T�A�o��a~��Vh�;�������Nq�/'�Z�7���'�*��e
�hŽ��e#1��bp%e(�B�ދ�V�Vz=C�J���T%�k�޾�+;E���t:vi;���_\��������LiU�����j�w��^q|�ݝ�֝}E�+�sI��o71@�$��Q��@|U��%�po�DE�Q�:�%���R�%�^A� �"���u���-M�ݘ��c��0<�k�����}��،��ŻO`��dJ�(@��'����dP�N�v�Y�^��oG;��*��b�7�o�Na�#u#syHhJ\,�P*��S���Y���Si4 �E	���B��fa����e�r�cf�I@���5��H�Ss��uy2�R��}�i��fK�Y�	����b9��7����}b#�ֽ�f!u-���}3BxδQ#���ր�Y+�����L0��h���	�>Z2�o�aH����U�G�S �,�ЁzO3,��!�wLIL����gNKg��q	��;��H�������ԝ���Ѧ��bo��g��^Y���Ș?NK��MwA�=2c��N�^n �����r+��V��&��Ͽ�.�ε ����T���C1�s�}���Z�v�؏�#��gzfٶ�ԍ�㞂��&�sCiQ���C �R.����	T�:��e+b��J����P�&�rTæ���d������8�Q��7�=�XZ�O����2�"��2J���.<rR;i�!�{�8��*|�O����ߘ`���:M��{�
y<�������]z�ζ��̳��H���m]�Vu��%���t��)���\W��������	:B.�����,&��C�[��%��~���7E�QA�Үh�"��Fo��U�m)J�>d��v�%��J$q[�,��֭,7�%q2��h��2Eȝ��Hj�-�:�a�SJ��fˀN�Lí�͒GZl]qa�e�������S��IỦ/�#����;�����R��@O�s#>�Z��V�ƀ�0��>����5��H�Z-{�a �J�3�{�y�8P�����o>��e��6|K�Cs�b�-�zH��\�d�9E;��+����i*S>���".X$t���pa'{�{h�`�D�\�[�,�̭�5���FN��d�R�B��oK]�9P}������z��us���&�TE�h}�k~r�LZq�γ����G�R���A�Iv
W
��%���9G�p��zv�/f�Y��1������u�\3�S<"h
��!�?��T�iul��B �T�{�	�m	f�׆��7#r�	a,Zc��g)]V�Y��N=��Tv�&o�c��NS�'A�3#g/���o�J)�d��SW
 Z�-����|���/��\i�ʏ\�jM��~�D�UAH
����@�ɤ.s�ܱ�ڐ�������}Y(����eN1��2��/��1Y����Y�04!M?�)��-H�c��>r����_$Ϳ�|�ē��o %c��m��Z� ����o�tO1�?��aބӔ�������r�?t%r�j�.-�O��5�A;x��(}T	Rgὶ=��D���\ͪ����D�o�n�?���ꝯ!}@�� ���Lmr���0��!mhf�^��na���%�c\�ȼ��jYQW�t;3HȃL�8E�KʡP�pJl�������o�^�Cy׋<��[�g�Ycq c
P�nw���"�I�� �np��t�'���`�m�'�~�oOfk_���/3��%a;2M��gih'.#�)���>I�$�)��l:�JԐ��>��$�C��u��#���aF��gL��X�sP��X¤m���i�� fN��W�f��>�k�x��D���!Һ2��1���+3�wv4k㎝h@d�=��à��w$�F�V�p�ޒES2"q��hP��g@����&�bfi�?����2i��	_��_�Nq+��\6j�kq�����mC��d`I��w�sM��^z��7
��}�zlx�b�9����?��й�!��o�z���Y��j���O�ބM�z���(*��^9��O�n
���<K 	���}��� ݑ�bm!m%��s<6ͅ nmqTL�~��Wx�oD+�)'7ɧ�P�Q4��.u���'.i�2@=:R�ۊ���4����X�9��;�E~�1�z��� 24`id:WB��r��K�p�?�	X�+ڽ��5	��+O���N�Q�_��	g�|��'�K���<S��4��Tq�v�� ��OE��m�8�0�"��簻����n!d�|儤:�N0�v�S���͊؋�]�B��8�3u�`4��{��������T�`�rH�Z�qzʲYv���f��\A�7m�f�V�w�nr��aO1��Ƶ���!���{�v��O��&�ŀ�1����{�I;�í)�`K��˿��w�ܼcEcc�e� �Y��Ч��1f̎�wU�*��-�3v�'�Qv0n� ��㮔����������Yᲅ�=+����CP��L#������i�oL��<��̈́�8~�qG��᢫�u-҅����˕S��|�(���b{�l��|�JW��c�r���C��V"C]��6@ռ�q��k�n���Y��͠��b8*D���|��f��T݇�lA��]|�qm�����A��J�|~n�y�6U�A^1��ϩ�"HŤ.�c�V<<d|C���&�X|�Z������?s��V����w,�=X~�>��d���g��{*RtK�H>;�mZ	2g�hu2UTiAjo�5X�oq��}������u����}%���Hֈh<��,���~'(�L_�"m��l�q0�G̏ &�7����f]�C4ˎ;���k���/�vr�.Yn��Kq�`�9�m���$�1�r�l��� ��M���#�v��R+nGa��^7'�P��-ԘhvA:{nL5��8��Wn��
r����" *<JT�!�@��psD+����<s�&�� &��zr<7G��4O���pi���Cؐg�D���ֆ��OfOD�:}��rº�pAĂ��i��*�r�0�2�
f�z�t�y(��VFm����c�����E�@���f����<L�q�[f�S�=Y5���0|�U�>�a�u�\8�0���*�x�dB��z¥���G��cS(sC��<�s(���'����6�h��A�!�w?�.�h݈�o{�YO���{ا��5D|.կ[g�m�U��ͭ鵯 =����A��1������J\Z!>M�-�/~�᪟PZb�d9����^a(�A�𲲮Ѐ?=�����Ҡ �iD���$�6�U�F��B�@�n�������ᄈ�\��<�Z@�u�&�A�#86'&�����I`(5C�h����������}�r���(_�1�yD۞��T�y��ؼS��Nn�$�3��m" Y����م?�.Vm�{M'd,�5,�!�o����~�RDe��~���(j0�ѿ��t�S_��DMt�	ð�rBI1� �u�6+��)VJf�8��*��_�� S�m��b�e����y1�y�}|%/S�e��G��|�Kg�K�<�6�bE+�T�����6����:WO����T�<�(M�FS��GFV�\�h�o�𥺢 տ,4��ɋ�@O��4%z�$F�$�ڈ�:Y���1�?TI�g���gBK���A��+W6�p�l��'���*��t��WL@Sx��э"�����b��$�<$��?x�X���|�^,�A�ӌ�qEx�ʪU�S�\%�/u6�378ц����l�ԺH���L�����}(�,��i��zٱN���$Qfj��/7�"V��j|۔��ڻ�����S�3
2ʊ#'�Wr�
��Rvg� ��R.-vk޴���A��B@RǄ�~���V�Ґ^0��F4�?�\o�b� v���)���[+���1F��Œ����d�fx9�	N�-9��%meՇb+����%Ն_���B��I8���7_Cg��՞�e+�N&��d�S وB��4 O��m�$����|Lj(C�؜��Rz����1�R�a���o�2D}����T�Eķ�� �5;�y<�O~"B%7��s�(
��F�����`�\�^'~<�eW`�,�C�?�-���b�g�>�e{��1����h(��K^u'�:��n�nq�����&�]�B?�G�DY���]x���~�5;�k�	F��3��A#����90O�,��<c ��5��R����"����C�LK���C,��G2�}�o�쌮"3^rY��e�"�L�af���{�U�򬣈����7��O���!F�p���}��g<1��~�**�$�<������=s��v�; [f�ym<p̫�=�{�P�aR�����G�n��NC'��S�.�c���*u�~��	�����i/��|I������a�g�i�q��3�,��e8Y|	��e$�#gT@�´���9K��m�Ks�<�3�xπ��[�A���u��������+d^��e��ƴ4�rl9^���6#�
:/�N8���]���N*M1K|(�cI�T��I�f��3���������)�x�H�w�+��\�h�^2S.��ZS=F�L�`��� �)嗜�=��9���[@�O�b����= ��@�� �[\@EB��
�\����P"����y<Of���9���׵: �N0���Cw�\���䉐�]vC��R���Ay��ڤ�E��5������޵� �S�������8W�A����u"[,�cTI��'O�wM�m�yE�^Q�H�JG�CK$m=����q�c3�˿�����h=�J%�&�[�WE��e�NYz�4�5щ����Z�$��4v-�N����+����FX��;�������L�r�Jm��,���	�С7�\8(C~g#��\:�(�r�Z��ܬ[����'ӓ�F;��^�R� K
�`�0��9�9�szm��*�$�w������| ��WǨ��p$�J��+�₤��s~�Q�G&�9:r���w�5X�Y�	զ��dvBg�B?��,�8�͸j]�y����.-���'�R���s�Y:�s�V�7?�c��	\��f�6h��N���J\))S��͖�F�-?�۾�  ���@�-��d��2������_܋/z���z�7L�Pc]0�m�{������"p������?�U{?X����rU;e�@?*[�;6��mS�V�Ѹ7?3f4�"�٪fE^y���Z�/GS�~���-��uɤ��4(mG�A&#��T��������F��㢏A�����cA��{|��&�~��a@7�N9�E�҈B�!=y����ݵn���X?�0��_�MnҸ.MO^@��L��ѻ����XZ�8m�H�mE1OL�'���id$�);���X����Х�'B1�3�N��8���f!.�m�k��8��l�ͱ��y�E)9��v���X,��yv�q"<E�PN?���M>[�^J�-��_��D�,��D���5z�F�	y�s�5:�ɨb�d�����v�	$�_S��	�,x������<�����s*�F՝i��-'��{\�џ�W��:�������Ω�^�,��k�C�}��/FS#�L��'?�I���x�d���>��c���&+�A�~�Hi~6iž'v:�����d�A�7y|y2_ﵨλC�0��X�K�b��ݿ����� �Ψ<*0!*RC�Ht��˰_�ܷ̮ ���ÌH%�}upm��7"���/��V·Z�l�p�P�,���γo���<�U8���
܍�̮^zV��(>	h\�>���ҙ�W�=��H��<u������M��;(N���w����5���E7�zy5 �Ul�l��k6��r �O���_�ħ�09�5k�`�H�C�w��ky�\߉�}ߒ�$S�5�vV�r}��a�eF��"~���s=|��q�gzO����V��巄���ץ�ȁ+���63h��|�K16pc!Rd�`�r���NԺ�6@5ͣ.�Z{�����R+�hAd��n�����PB���,��Qa$�#<e|K��u�DVh"�g�8�AC���IQv�9�*(�����i"{�� 8��5�� c�r6D�
�W�w<o5�P���{�&6�v���g�R
�ƈ��Y,{;&��"�l_n�O8�3?�b8,bj��Yњlr�1O��b�Qd��:t��� �a��_\09,<̫LI�jv~U�Еǁ)�V�sP�'Jw=�h��%���i��馩�g�%�s��;tE�1�J�Вs���Ș��T2"	�ej*I��o�4 (���$#���F��ʓ
|2�m�mm#	��lB�粢:�v\����u��'h�V����V��GƜ{�� �����^�ͦe^�Yׇ4�y����Y���L��i���c_�,-�[Iણ�����H�Nk�`�s�勉~�VN�U�G;Im��m;�m����:��wh��A6�����Fh�,qۨ:��w��F6�d�D��=\����$G�/o���ŧ�M�1��L���c���R�����`\��Qd��sNl������d6,;Ɗ�S�D��L��RB�wE;���J���o3�` R��m�b�b��4�b�BK�7x�Ŀ�3LY[H��	2���#�Ae}A
�/R|
�0��5��R�n�N���R~:ݲ���GV[���|&����f��ȩP����[{,n����aR,������o���43;5� ڀ�O�	�F��G�['�F��J��q����� z[k�V0h�=OY4���J0� 	���󆘕�		���2�'K�s� �G�,v��B��/:��Zʲ$>@��?:I���L4#zo�u���K��5	���8ܹ2`�P���a��)2�8@L�kg�	�nTF�|�M�E��qه�P� R�oj�&	����� A����6�@�w泙���(�a�$�G@������I�Jb!�Y�,���+�WYk0`||u�G�T�&Xyœ4���2dFp�U�I���*�4�ֹ���WeJ�y��N8@G��[�W��U�0[|sN�F]�k0�q���N5�����tO���r��QZt ٞ@�pn0Q�O��-��:�|ZVl�Ufy&��W@S����B��t^�]q�q�S�3�����<�!P���@q�3q��iq �A��#�0��uΗ��X�|�Ǽ�D�5�<�> �ĳ�O�#B�B�mv{a�ќ���2N�����	ť"��EZ'�|-���D,�r�\��l4j�Ԫ��I|󨘿i���nӐʨ�v1�G�l`��5F�L��y'��>��u��ẘ��-�PmB�|R85kS�5X=`�R�&;$%)��~z)��m�@'��N��d=C�.�M��2 ���%y�z������� �Rf��yea��+�3�=�h^���TՈ �0����:.M~!!���,"��-��Smϥ]�C��8�����-�R�ȿ���>DG��/C����G�}�89��+aDY��/!�1� a8Iˌ��u��
��F��1+WI��crW�����
��(ܴ"����.�Ib�m��|�O٦O�L\Bx��J_-eDN��Y�ú�xa>���M2��QD���5�$C��/��HZn,)̈́�B�gh��^%��z��f���ڍ����8~<ϝ��@�[������Eѳ�*0ز���)\���.l�}Z��J8�,��?����%X���ѭy�:��"l�=G�*�ٞr5���]�^G�6H�P�,P'����'ލ�p���#��JN@���Ck$�&�����p\�$�bhi����(��Y��O��`�F�Η������F���|_�O����Y�y�w������r%9e�z���vj���ȣ���"�]�����AN߲�Tu K��c9�!��٥p5��<*7z�J�-D��6k���"�M�;Ws8�S�j��6b���[ M�nC	^�_EN����V����*��˸�{(#���)��6�+�;�,�{*�́-��<佬v��3���s��̰�b�|�6�����?<����a�Vg�[�y��!�;){N*p���� MF���!fv�H����Liu7z4�8 ��@W-~�w�:l���&�r9��3@�����LDI����x�]s�%dre�
 ��b���6�`�#v����`��- �'�CcBe�ތ�K&�9�T6�*���_U��L�N��FY�������}@������m®��-r"��Ļ����y���E -�_2#���u��h)�Aw	���,ռ�������Le	�x3�l%wB���?)�;���c,{D�LB�''j�$��e�WE��_0��=S2�A��D�$/�Ǿ����9~�t��M��tdtzJY��f^¥BIS��M��1D�0E�#O:��nZ
�}�SE�vP��_$��{�B��<i"(�R���*!@��͉2\]��g�W����������z�ې�{k�i1�sU�FR]o4j�Kj>��h��9n_��`|s���2���!�g��X���XG1��F��l��!-R6Ff���mn�Nl$�T�E�R|�qع����8�zs���ry��V���*�O�l�����8�R������{pT���W~NV��{ǱVԑ���՞�1�����Q䤡�/�.=�(V+@t���0��Pdl:*�h���=���ڍ^��7X�����o������N�ȹlۏǶ�.��!=�g^���<��}�evlt�h�9;��������X�N�[�[ǻ�}qBYM>\�0;L�.Ik�K^DF�|�U$3p��G�>�2zl���sVE�K�c+�aX���(t�*�9�`7���pS:��M�R���W�f�)�V���.O;w�2i{�'`:ʮy��t�|��i�:�!F�28w���l3@	��١Y;���
�'��i`V{����(�}q��k���#�n'faG[FaҘ�U0h�)��h���Wr�h�I�������=
��2:����[eN�c��{"�A6��uq�I#
��S���y�� �Rg��B��G

�[YV�%N7�U�G+"NwB�ܔ|�E�()���F��p�-�d�UhP�*� \r/ q~����������|��uq��8��E�5jՂ�b���>���&�zGr�� �8��S��/Ʊ5jg�dA�.��Gq�h<.����@��H�Ew�=�'6b��#sl0��+}O�nHq\L�O����C�G��F�<�s��yS�	R>2!�ʯ��ú���[-�֦:q�z�Z�Dmz�F��j��G6����s���J%_�#������w�}�Q��y�+�6��G�w�s�S!��ڳG�`Jl��\����	����:��L�YK��~�h�T���0)�OHH������O	��^'	.L)B[kw�먥�#�3u6�;4�mB��kܜ����4s�>B���P���l�	���O��;�"~�����,��/����A�W"�r	ik޿ՅW���L=�e!s�38Y���Q������e�O]Sv4i�;^x������8��z�z��r���ғ�®��!I^5�\0��G�1��)<\;���>6��vͷek"��i&I`�SG�m���o��Ʈ�@��}T!�zb�iSf<-��% ī��p�8��T����[�&�:r��;H|}"��pn=� �q7�� �j*~��=w+Dt/�C��=���]��D?��#���F�v*?��Z]�����YH��5*��L���{$%��;�%��[u���W��-b��~
SZ~\]�I
cS9Ϟ�����<�?z$�����S���b�z���_��O�ø�h�8P|"���Q����m�h�/��!9�A�n�>~�����m�+G�bYY^+��a�#h���e(%n�-��9��.Masn���!ʹ�ӕ�N,���6���G��4Ea'�9���.�4�2�+~8���I�=i1��.���`�ӂ/�A�1Q��H���|}Hq� �S�RXbc"�
sK���h��V�e<j9m�Mn+���H��@���>*�:�\5ߟ��~;���a�au�G��=�;gH�?��. e~������T9��x���R��"bF��b��0Q�dt��:�QP��L�&��WD�O8������w-�5�v�Kax� ��<H����fx�"l���h<}���@��(%��~�	�� p���xV�}D�3�����]��\v�
;�)�l!1�7R=r[�V۩�WY��-�v��0J4��A�@U~���0%O��}z���_�b������櫖a<�3
��K�%�|���p��^K��E����/1�ƙ���uH��=�.3�楉�ǡ	���։�T��֓yI8�aZp�V�ʶ��J��eB�KM���q����e��v���ˇz���^?"�h����=���<n2N d��ʣC/�)<�SE`<�IEG8]Q��ù���Bz'�%7K37@�،�5�v�������H��K��o�<�3�ܞ���τo7x_�'�+�h��N�� ��Kd����p�DlP��'$g�#�9W�+(7\M��5Q=��c�q�:[s�J��T�p�����I�@�3�
~OVh1��c���	[0<��l�3k.!�B�'q���T�hg#~���3�S���	Sb-��D�-�~Ci�> )����T�vm'�U��'�i�i��5���Ѐ[�X��?�]����O����R�M�͹w��X�k#�p�O�)��9I��f6@3�����l��#���9(U,s4oF���{�t]hz�@,���O?��E�	�`7�9��OͳF{�Dj�R�uT_���k��B�𽾆��#	�y@�J��c^�k���¡�A����1>�I��m��S�w���)bރξ Mg�{i'�������"�sg)&�����sE�hZ��T��e�fD+ҟ9�}O��[]
7�<׍{ӣ�b���WL�x�1k�"���ՂzMAƮ��t�G�j	"%p�}�%7Xa!�>9��$R�p�B��h��oT�$p����bw-��:��Z� ��!�[\���qvLY�uM�cb#���eu�M�tf��a�G(��0�e�qg�2�8�|"�d��7�	�qz-2���۠��ҼT�-ְ�ze�<��{�pڋ�S&bƥ�"�������8p����&��t�U�E'��:�����J+0�>�ց��2��2f�/U��0�$��hRĔ�6	�-+;k��/�M�kvt�~��8�d -8G�y�}������뤬9ZsJ�����ѝRmEHl2��[}f�����þ�GI���)L����\~0-����gh�+����Y�X���GRR����<֖��G��צ�V#�����S���vS�z��jY�|DaS�˜�����!�������T���&�&���%��#U��֌^*�Ь�# y�Ց�d���½��7�LiEw{P_��@�lR3� kWt)����^Gc�Kj� Bo��>�ݶ���fA� �UD�Bl:�=�p ����~�ata*03��*XV
��
5C$F��ū�Ạ'�y�ȼ�l�+����b�~��M�>�o(��&���=�l9�B�2G+�0� �ޱ��Čd�(?@�]���M����V~�y	b�l�0lwnZw��N��'�#֥:��$��ڿ�h���5�fp�q�f��Q�Nwg�}ON���R��B"�^��gC¶l��	^+�WǓ��\����R�kKI�����{�_�	������d
f+-�F�ō.���;)M$(����ӷ�q�뿐���kD��jLz�}=��Ӹ��}��b|YD��l��`�/s�xj�=�xR+C�⃱l��_Lŝf���υ"�����2W�Zk����&3y`�1sB������:׃",��������ʟQ��[:��5���e�N�t��D��Y5�a��I-:A���z�C{���4��o�@���E�=V⩔;��ߧ<껭����B6�{ac�j�ƢIz�H�x(���B���ݻ�^��k"2b�ኵ����Wd<����/���"!��3�o�W �mPL��pr��4���eg ��;Uh��B����JǇ�H;V�p4}�"�%�w�hO{]�`�� ����e��cW3f�n4;��!����ن1��7>)�-��LOsxu���%0��7�4�b��d���>��#��M6u$����B7tRlq�]�φ'~�m<��%'o�d��~�@��by��7t�aoV�S��z�_�X-�p��_7E��.\2���"��usF ��s��I�P)<��[K��1�Jz~��W�Y������X�>�� \ë���/������S4��&��hT(=wN֖LVZ�X��S��V���6jC�iE�%�"�oW�lH�ū�l��_hcN
���?[�wQ��]��h|cwQ��CS�ꞹ� 7u���M�+sOWm�!7�{W���}���.#�bZ�Tz{�dDc��w<���t��x��&$��%w�%���^Z?{�3�,�
:��-և�]D(�!.h��Ѯ���ՈG"J@��0��ֶV7�P}��ki89f�����d�Q�sa\�ݧ�WP����S��~���a�H{�]L��H���c�Bt�L�!�6E�jE���NbDwB|�Y#�"V��%p������"�� !
�FDqT�^W´B�������O~��n~g���D�0����vn�2ڸ3�������\<�D�+�g>ju���;TK@jE��j0|��놄V����E^@��>@�UH�3���%co��~��/�C��R��Zg���$i��N[&_�lS����Tq���a�����J_ ��bh��[�!�d��<�y7~������#�n�@��7`˽Ě��&w���H�9�Ʈ��~0?E����*�3����N�z/�ќ?2���t�@���ckP�`�Tן9�R?䥬�h�y�'��Pri�	7����/>;z��h�_���<�z�t�;���+
���z���}�9g�B3G�ȬK͉�j��0ߛI hcbqY���ό~#�e֠N&�Iv��<��'4�=�_���>���X`R��rC�J���Vzn�n.=9e`}e0ÜP�d���yL���C���5T���9տ���y#�uG�r5�ܯH�ޜ�(��[5"ƨ��U����������������~���vL����.ЅD��7���ȴ(3ʮ�n����2����P7�?w���E�_X�[Aa`�� hpTR� ��	�ѣ�%BV"���Ф�XZ����N�ē<c+d����E! a���Ր��[P/i��f�h�5;2�.g�����"7\>[l��~�f�����9px"t��Y�x��¿�q��RT,c�W6�Q��j/����.8� �mv��+�� ����`>�M�yKp\���A}^t$C�Kk��Ci-�1�XԈ���[�BUK�W���a�Z���תeU��4�(�Bz�����o���f�5	j��<K7�Y�X4���~���hB�[��')�������O�;�2��[��o�:wp�췿�eZ�V��# L�09\�o3wy�/Ħ�BAsl��}$�g�i��r�Y� !���PA�6�W���qI�ơS�Zb{q�*�M�Lf�
N|uq]#}�͙�7>�B%�{�{P�O(N�x~�����d��k�CbzGut!ji�.DE�k�QDl�`�t�26ŭpM�V�N�8���[l���K���:-��y�|w���w5��6}W��5_�e����#�0�@u������(�j��8PB�􃸥$��?hQ��´�;_h�]�e�KV
8��U��47�h)��[c�u#4�d�}EpY�z�~_��яB��%#�-����́��ܶ�9�d-/RTg���=U�fOR���_����gs���,>+��nd���5b������PaM ��Y�.Kg:ģ�e�~��̓���_�y��(���qz��v^�lC�u��H�E�@p
���6��PE��k�����;<ʁDӮ��E����H���?�l/��gˊR�t4q�΢5P��{:�˚��
Ԥ{�r�=f�UsJy�!�tPƼqھ��Hls.k~F��ǜ����g4�E|ʨ��_"ͮ����'��xuj,h��_�N�(WcF��u���y�k���v��)i��A�?�
�ތ�П����Ma԰I^}MG�n�8���r|M��i�ۚd�{�C�F���F=������#B����G�e�h�]��é� �s���x��x �S�IHOzR[�^Pwu��ҙ�i��3�N���k\�7b�R.7����ݤ]P�����7l�`
t_^�{�~�N�q{/�a���3�9��5�"�ٻ�����wԁ�V�]4�/&�w|k���'�A�&�yb��CY`6',�s�U�m�g������S�����&�
��n.��s��4�o�����٩RX�ӇR�+*Qn������%�+��֞^�C�F،�b���	�Qh�y�*��#�>�/Q�~�Ou�������B�L9�1H�HK*ZW��Y�"�խ�V���"�;{��T�e�z�5���M,���t� ]1��uKH�I�n��ʺ,V��h�b��U�ai��|���C�.O�p����:�o����s�<hK
�f`OX�0��55�h����Z�:�0f?��G����D(�fxQ0�����ҦH�PN��s��5��9��=Y�L+�����"^@"Lk'n����Vw0�o��B>PR���ٞX�u����	o��ԛ��Xİ���lLQ��*�
|1�<���BA��"�g{�M�$}q3w�������%Hy�P�"I���F/�n���Me#3�6�o1���~9LP�O>��Pwa`��y��~ǕU8;-�c6$b�S�I��wc�{��R�!w)�r�?I�һ:#�B�D>����Q��%�8;�mX���6u��e�J׆��&5�EP��+�����/�jo�)+��ʰ�0�K�ZȦ��,L��<�xchQ��MXy�>���Su��#%�<&v��=�����/c�J)ʂV%�z��gH'+���v�6�ʦ�y�HB]�! �*��)�N浿�FK�ĝ�S@3�;ʫ3c[�5���_� �X%^��x��T� �{d���m$�X�U�Q�Xd��w��/����
8�@��cɡ-<�Ƀ��֜Ǯ��ia&�y�q��|�"}R?�mq��Y>�J�u	����	Wj��o�j�/	6j�Dı��l��2��˲CA���r�b�Й��r���O:f��:D�Ȩzu���J&`��7�v9`ך^q6s$��'����ʻC�/�dvC�(��&_��ǅ����P���z�޽���8�|�xx��bR�������U�6щ:f�|����+\t�[�3J� �Uj|�`��OT�k.��x�����m(�@�p*�.>J�{O)r��H�i��ݧ�A�eHg�g�^��+�d�g�;��% Y���eǌ"^ȘjC�{���p��I������z8ʪ�^��#at�?ݩ]��׬҈W�`���ᗸ6�ˎ�HU��J=�.�0,�ay_���~q�q
|��$��0��Y�wK�l2�)V�LC,lM�W��?�x�0��OnR�&Un���!/P�:�gT��%�$xW��<���`)+��~f	k��ݧ�@a�����)�v���R0�6
��[dx�I�<YMt��9�O��I��� N`$2l�*�l<à�����Q)�&�ףO[�*�/�r� Oݤ�^��X'T.����^�A ���=鿟��;6�����RwbFgO���hK,4a�p�JL�82,� e��l6�� *�(,o=�_��*��HB��5����FX��O�Le(�@�_�j�o�kSȧ&�k��ں48W��֯����tW����T�
��Q�sO�b��[On��2�������/�:�z�N6y��܁�@x+�F!n,C��}����x�K�Ԇv�,��{������n�B?��$�:њ0&�n�Z�o��S>�<�4� ��h>+��5��GmC/�#�y$To���l\��C|=5(�8!�v7$iY8@�}�{;�X����F�q(A�ra]/�Jl��k�(��oV�<P:���?oBD��0u�i�+�+bth�.��:m�ݶ*�	�@��
�uTf�JV<���$gI&ְU�΢>�Ԁ����H�q���un���m}:k���͍Lt�{F_�~������V�B��w�:��G�|"l<>��.��ӚU��D��`(��ӿ(��/}@^�^���U�^;����S@�s%��cdOud����F����L,�#�\����+�g����逽r0m������T���%�\93�Mb*)�����4����b���u�F+W�:6���OJ�|��/ IϡL�C�~`��7 ��67J�*�A�(pE���[�I�G\��g�i7�c�S����Gkx҅1M~�oY���I��}�A������/��1���aw)`�����K�8 {���v���˺^P!W���j���/0��.� �-��G�T�b�	Ҳ�F-�����{�����A�(�;	v�'&.�sdR�{I3*�a� x�=��aNWɉ�)�D��3��;���Q蛠J�%6k��{�M���L��@�^��
��r���;Rlq��jk�a]�klo"-���lQ�,��/�#N�q'�t#5�gߡ��o����Ы�Y!����"N Ȭ�p.�!��W�2�K#bD�&=
ȑn���R�NQ2x��o�GK�zKv靥����X��PeN���Sl�b+U�o2�1Q�/�v���6H�s��>�W�д�F�,C�7�w-�#uYX��z>���Th{Y[ta,nn����TqGfV&+��v���^a�j�f�w-��'\��m�
��6'
�"��癛H*q�$��p�����������Al0��,,��� w�u��2]�_�Oqvmu���y��u�C]熻�WQre���O��U���
WQ�oN�u�Q)Hu*�� "jNeq��J�kn�p@��S�xZL?u���s2��\4��f���~���w�����n�6�¶�U���B2U�%w���z�,��ݱKi�l�t;����7x�*�&��<��(`�lF%�M�� �h;�(���I��&��
���J���[���1�9��c�ImIS��zW�u��N�'��8�
 y�ƺ��r2������(��[�� 8K��Q�eOAx<��5�t�/	���FaXe_n:ͭ�sH��v�ZЎ"��١�G=Ͱ�8� ���bΟ2������g)�,�8���}��9Q�j|�Ԑ����cIT���S��y�����pq�uA��Ǧ[gϷ�t
�V{g�V����fGs#}�r�T��2F���`�=�W�T��1���\QY�g�=��VD���T�a=4���J&5��Q�� E=V�0_l��6�{��<P��#E7ЉV��)�ݭT� x���_y7�X$�s4:A��,�ɥ�5����[���}�g-0麹��HO�Q.��؍�5�v���גک
��"�Ԅ�ξ���t��=���J��0����z�N�ǆac:U]�ɣ�SLEpE�ܱ������|�u_k�0v�����Ĉ	G��2\ �������)z�}6sR*X*�p9�-�8��s;���lֽ�)�`�[ճ�.����������2�uZ�1+ D%�9��VPQ�����9���������6*c����sTk\mБ���2�kI�~h�@�UQ�7�B/q�-f�7Eg��a����|'�ҷ��sP�4Y(��� �N���G*�ѽ�x�����C�%��'�*<s}|O�ؐ�<f�[��hu8�#&2
�	.��(6f^X��^�ټ�g������w{x�	��/������Sj"e3$���j%Z�����&�9�����ر&����2��AH��OS��I�Z��e��v���<U߬k&�f����-Y��(�LU�ۃa�^���+�gP X[?�Em`mS�f{Z�a��3%o6AS���N�����xh���vr���G$\�E�ޘ����GB�w<��A�L�Ԣ��� ,`�&���3��㋛I��2�ߣ����eu�Q;@���UF��^�'�2bW���� �H|P�EDݚ�@b�l��K�0G�r�3��y_YG�� �y�$���7�c��`v�<M|������ ���4��r��=Ò�7yϩQ%�.�5ž$�#Z���FK��
�c x�,[-��u4G�Rk�}��f2H�I��o��?�ⶢ�D�����$\��(لr̙�WN�&�x �Os ��*��&�_�C;@g��!m��L��L����}��>��,�je߿�:\��M��#�V0ŏ�L���!��(Ns�e0�׽ �LR��M���
�z���=>��>�'x��F�����i	L�!+����qMݘ����dm����hC���=����%x�*�<��&�ai���w3�l¥U�#rw��5^\�ұH=��!�(�dio��G_��o��t�~cz�u?���D���
���=�����
,�w�r�1�n��D"R�&{�1���8�S���U�L�#t�C~P�%��X��.�dhoQ��.�C�B����Q���As�ӇV�>�D��4i�뇰��Ic�`i��a�=EX��J�!�E�N���lx�����#/7�F�|jI!�%さ?��8�yͤ�(u�ѱP'$���O�S7l��?�qls4�'[��$���A�2�T�?r^��MƁ�)T�p�wD�.��;(]�Ww~���d��h�JQ�L�{hW7���l��,�D�x����~!?6A��C�W��ת�P�ېc^���&�t�6(��ފ��X��4v��d� �J27�+W�jEu���e�Tl{7Q��*����,/a[/�a|0?I�23�S��]��R]�7ڒ����ᒳ}z��.��ӆ�)���v[�ʋzw�5�~)�ƂP���jr>��7u��HG1P�G�j
����	�U���I���.+���]�+�|�AR�)��}�U�i���R�����['K\ոWu�u��Q��������sq���X�J� ��a�Cƻ��J,�kْm)��m����0%�9��7�tɧE��n7F���#�@'Uр��M\e�՝�����I�GMo}�<���b����O^}�f�t �_�o:����D$B���l��LER����J\rgoE=O�'?�+*^����"��-�P ���xX���Z�]]���*���FD8G��K_�-��m�`y�Ö�S{�&0;]�<Q�wQ�"�#M���+��esZ�%m�5ܲa��YOW���T�}9�?��_�?(��1�x�x��]��[���'��wC{����[�
:k	u�J���Ƈ��7���8h����-xP27��U��ɶ�A�/�e�������,���]n|ǩ�d�+�w����?o���n� 4A �O�Л.���|H��1������n���L����0Hr�!=T.�����[�%�%@��bO~��D�Nt
WC�/��&�y���*|��dX��vJ,�i`R�Id����u.�|SM��F�\�e�`:�@ ��f ��z�1	��]�/��5�T,�,��ծ���������>Yz�zA^|�Jk�������GVܑ+9����	��HN*����o��+	�^��b|6�ۼ]�0~�2&�	SnCIs�}Q�@�>C���ܝ薣I������,u灀����F���Y���y�������z2�R�(����pk�)|���$�(�Oj��4�Xx����`�3-��])�x���@$b9v����f�%��V��ӆD�^˴uz�1y������,P��MF�J
09퍓�պ���񛓱�B"2�'z���W���Te�@��\��
�bs�e1u�=�w�S�71����R۰:�N6l�(��𖘸
��_�~�0��S��#�̽��G�ލ���[`
�_:�뭑Q	|�!	����[e60?:�N1]��SC�#/=
>�.�I�$����&ŜR]��������F�}��
�z��Q��ע���ΉF�؁ө,�&��C����nq�i��z"�x	4�3����r�:�:��[\��5%��_��?��+ ��Y��x3׿�avR�,D���τ+p:����)9�������dc(��+9�g��C�N@�%:�<j�%��#��'��� ,	MP�;}�>���������r3AT�u� ,h�n5�]�F�l�'>l [�9SW�1_n��^�&���${-�Ͱ(�!�^��*@8�z��R�pwwrN�dG}O�7#`�6��G�jC�~R�r��#�*>�2ג[�?���<���g|�~4��ǭ��"�R��b���m������:I����7⌅ �ZֶD��rV0�hCg��h�9���^T�r:B�����Uho"����{�W�y�\�;�D�O��A����d�2�c��^p�5��u ��\!g=6 ��(9U�:{��i �����]~D�W�m��̄S��m�7UI�P�@�������#T��*��
	����.����@�� }��
p����u��MY]�e��xn�N���E-q|Ő�vZ蓆1���,F�^�b^,x��'��w�kϽ�������@��@�����#W���(��H����؅�ES2���M&+?�H���yAy�Z(��i��!z�7���7�t��֕S�t�e����*���`����r!5z�-��ԇ{������|�Z 
{��db�����y\���%�\j�&�P��Q�Q<!M�����y[\�����2粓��C��d��GS��q+rz�S	0���ꂘ�ŧY��~	%R���j� �O�4l;-PS�jݜ�}Q�kb��:����*��m
����� ��Kf�_:U���U��/Z1o�&���KJ�D�	�5<�My_*G�C��8����1�B�d�y�v	P��g]�Ŏ�/h4�"�9��u)^�{E�Cp�>�7�����e��9� ��P|{VN���)�� gJ�
�Y�g�[�ұ�"� ͂�hS�ݵ�5: ^_҇��x��N~�7Y���ed
����[&�����	�7�*C+�Mّ;+��KKʌ����(u�m,t��5�\4-}o�����[1���oyvN�|�gh�d�w�Rx81e}Y@���o��ڎ��������"xpK��QurÙG�"��� _��ɿS%i>���QxyF{X>���]��܄���~?1UJ�و#��]�w��v���]�R@%� �Y��#;[D����ܺ�
Ζ(N�}_��cW�D'���7��]}E�}���8:��I�-�u��ߔ��E�6�"�9Q�����z(r{@*8+�0��{�I%����6�4<,]��Pp~���jD��ł [�;�B�qWd��ͧ3�ۙ{�{<uY�\N��pV.����L��͋�8��<݇��}k�{]�&Hک�����м�4��q;�Av�d���p�I���"RMZ�#����UQ.V������/{s`��W`!H������WgIK̂Wa�עȵQHūEז�� ���� ,o�x��p�d-����]0�4�+�&��E�ܘ��e39z��L���=-�S���1�1W�~){C�������0�gE����p1���p|�P��n�����鍧zo?S���@
〷������o?��c"��l(惇�J�O��o�*�N}h+�]�/�7��#��H��A�1.w<��?t>w:�U�f��z����>���:gؤY��4g�}\�oPШF���;��m�0��
���J#X1�e3FB�/��õJu�����7��H���[�Z�H���UAm�>�5��˓xfv=v�3
�X�2��ލm����]������8 ��:~����	ȸ�Z���C�	�*����K#�ϴ;ߑ��+%��=A"�lƍ$��Uq>(��°�㜧<���xb�/����E��b�A�����~�ƪ�R�7J��<]3��bM���]	e���-��?+;ssF�����L��/m���;z�4�2Y�
a����n/u��r�o06��E�2O�}�n�����5h5��ZyEY���K��{��`��q��r蝼j���n �U���Z���+B �GS1>;�_t`��/�X������h���r �A���`����?�۫�פ�3����z�p��`={�44��N�V+,�M"_z� h��z0�����p�}�O�]|[�[Pe��9�A���^5:Ȫe4:^�@�D"���g�3�&���J���J@k�,k<��v��V��w�ݽ|ß�����g�P����haȋ�{\g�n�,�12�쐹� c��Z�r��]O�,��O_V<��1�kzސ���I��UŅ���
�8���RyJ���j�-���A���ҔA�d�2�ܤ�[�5��^�v|�nW����Y��|ԇ��3�v�f��,v�E��j|��c}��燞��T������68��Nύ	
�7I굫�*:q�]�bX{�P�|*#�(��	�c���T!� k�]?[��=p#�ʀ�-I=^
O��K̖`s��N�'�H;�@X.�}Q�X�D%�c͕h��G�q��L�>��S�9Yj��޽�V��.���U��z-vN�K�*<��ֈ�����S�nؑ'$!��3˘�#�_~��^��| ��NpZ� ����&gJB��s����)ހ�
-\�A���m�$|�=pI��R��j�(l�J �;�� �G����
�Z���d��4�4O��
�'�(����/�K��*j����/ʫ���II����d�Yz�u#�,;A��o�3~��ن�,υ���w���dh�w�Xpe#`Sv���>�<�g���lC�A�)�j��N>'�i�d<yl �@eg�����3\��vl�j��(�b�xi�	�3����~k��H')�\�V�f�Q*T9<M�XHqE۳�Ue	.=?f>o0W����+Q�b���i&�N�y�$:{!�ӂ ������N�kκZ�`����~�;A�ߺ�Zuj^ҙ�Ļ(��x{�_'+B�)�,;z���j���Q=}�/,Bs ��.��.j��U�dZ=d˂��8P"8����H1ݼ){|�u���4߳ݫR�,f�����y#�o����E�Q�e�rQvD�nU�Y�;�e3uJ,����>	3�����'����!�S�vD�V��xZ~d���!�FrQc�(J���e]D�:�/��o�a>�J8�һ@J1i�:SI�"C��d�|z./�wٕ�K휋=�Zy��gslqʄjI�~*[2WjO=��p/��wQ�U��]�-����okcp�����Q���_�AB�;Z�kNg��9$/vU�v�Pr�(;�k�]z�i-��yFr��L}?H��T�yՄ��6b�*K6Yh$�B��5�ް)¿���.8!�ڗ
CZ�R���ef��+F�n~Ĺ��nn�(��a���"-��D�<�	�4Ԃ�ݕ��8�43	H� ""ݷ�p����c�+���@�Oy�� �)�ð�ԟ�� ��N9���(����ǔ=��w:en���rJ�I�y��zY��I�4�ٸ��ohY3����Jq{'�F�����N���w��5G��u�M��ҤO�4��A�I�������!�y��*��n-,+}�L0Y;')}<��̟��H��3�����Lo?}ʺ2VS��z���-�V´��|6�o���G�k��Wպ(���K�޿{�I_�)ף��R+2�����z��~o�K��Nf�I&<f<��^��$NcR����8���8q����+�����S�2iRU��Z@D��>R�ʆEX2�d���&��Dj%�#�@�dwR)�ծtE�� �,_O���M��(�/m1�H�� �����l�����Aȳ��n����=��+`|�x����l��:rg��	���ᰜ���I��!1~�S��{�"�x����\�I� �[̉��h1���u�g�^�|���������}*H��k��  �q����2���t�b0��7	U�.2����	&��� YCX��)c8�grI���·�~���Zz�D��Ţ�J�� ����8��G�f�N�/U������u��g�ܔJ�L��_�(DոPwR��Q�R�W��#)��>J�0*�h~v��.�u�]����V�Xb��Ѥ�-LM�*3�/f�9����ٳ�1SDi���X8����j��r�\�6|����f�/R�im؟��y ���iO詯.�Ԃ�Y�S��,�L��}}�%�;t��9�Oz|���u�[�0 �(;���y����a�bV���	�mC����3pz++2��vA��f�<�G����Ğ��s2�[p~0u�G�Kz�A�^�p�� ���8��	��K�-�i \�W��%�����������
�mh	ǰd7A]	�u�����t�r{M�5�����5r�����u+���:-���A�T�z 8�re,/���)q��Dɷی��أ��ړ=���Cz� �t_�����ln�/[h�I�TY�;�/��p�q��bDQ9�#��/!{�1}�6u-|����/C�(���ü}��ӠU�k>I͈�~��U�L�xU`���K��z]�6���@-#�XE4&��F�{М�)�0H0��u&#�#�h�g�����i�dSJ+hjby�`Q�ebT��I���T���:Mm��8~�M���d���D��p��R��>fj�T�������k��yoYI?�$=�k�R���_�Y(W�񴹧��R�?��iw)H6C�H\[���tq-$20��!��9;�%�d��j�"ԉ=�;ʉP�e#��a�d��i���܃�#-4�-���K����y��G&�fՓ.���;��/_���6�@4,MP	�zW�?� <��M]���b�Ԯ�V�,�f�}U�G�y�Z
#��wb���L�Hd3d��]�Ñ��(ef����5w���_�sHb��?����~��#�1���Y(
�V�0��1eF���}f��v��jP�p�/*ND W#^�d�$���w���_fB����Hk{T�p���3t��G K�G�P�	�5��dq�0����Q��~�_���-Ͷ��~ڹ������<�n��&i��?N��P�u�ʻ�R����N`B��ZK����31u�Ԫ��D,&�㷙��b!u��.}٫���FD,t�h����;{��I��#�^�̈́�W��1iw]_0������:�AD�1��U"W�].#}���QA��j�3�|��r+����A�iuʳ�[@�ͨI�ɋ�7^qf�<=��W5��Z��ʕ�A�X��pj~�w(�����q�b����aɘ���l�k$�Cp>���%J���@���`r�?�؍�4<���.{k�=����{,��ڹ[�{�%�������!y�<E}B���t�2��8��E�Pep��$&��M_�����.`��a�iΉ���������hk۟�@␎x�TmS�<S�9�ˑJ�ȑ����[��G�>Ǽ|�j�����Cr�����"(�Df�b�Vu�[��������Oϛ��դ3s��?�w�Xz+�7`_�hm�PwR_�
!�s�Ѵ߀l=́�K����kO���E�$�ϙ��kw�4�9��U�������p���H��t�� �����oX�E���]pLW�Ɏ�,� �dߴ�%�3���р6hX�>ᴋ&��c�}>�Б����J{v���(U��>���S�,�!�2���h�����2QViM����2�M�}�C���aMr��J���Yp�Yo��<)��bl~JQ��_�Ub7NM�S��m��#c9��K'�>W��;T�#:��_�^s8����L8��}v�Aߏ[��g�{s8F g`��1��~hA��*Q ��w֡���S��}�n�΂ʆz�����M���Ҭ<�X<��zr�p�!!���i�Ui�IU�A��h:�=~H�q#=ĲR��t�<���y4Nk�Vl7�@��Ⱦ� j�睇5�غ�e���������������.�j�+t���k����k'p�\TE;�33c8͍�:���A%1sFF�\ۡ^���U���=��7Pg�w�x�*�/q�w8�X�P98D�c��&�8�rr���x�6D�Cj�v销�����Zo!��"+��h�Ci�i��U�W����1Uc���rRĂ@�	��C�ۑK��d�;�����2d�d7@���έ����5�B�P��}�!r�n�@aA�g��2�C�~s�_g��4�o���QޫY�'f!*L���Ӹ�ͼ�L��S+O���7�Չl�'��GY�Y8�̜�Ɨ����*�ϸ/*
��K/9>�>3�g:6UK�N̺��L�ĉ��9-�g��b����V�ѝѐXm����48�bO1��ڤ�~{Tj������ב�(��%��F��b���4� _$N��6�]��|u�J��?��iuT�;���Eyt�L������֚Ӈ�~��x@~h_C��:��#���L�SMa��r�[P"vO���~iw���>��(��c'*ף�ȷ�g�C�f%�����p!�����ثc_,�6�3��3��d���9����K ocs�xM ���!�\�V{~$&�g�p黎Kw�Ov��)����-\��$����$�q�!W�y�`!��6�%@�1)�ѝV��?�V{���i�fƉ��O��$���أ_QŲ�"}@ߡ�5�����c�cX��	�K^Uݹ6���M��Ek �b�e��/-m�"T~���N�z+�z�d�Us��A����a�Z��UpF�]ѵ����-�ږM�����Om�1�'�ɂ����Ύ�j������Q�ޥ��c�ȢSUMI��f���+e��^��rG�|6����kb�ͅ���W͍
Q��z2P4�2j#ۡ���;TBἠ�X�S<̡\��!��>2����$�T�NQ�
�M�7���V%i׼����'����ވ/�R�ٕa��DLY��fS�/�.�7�%_y[;X�m�D��>�o=�Dj.Aa�rfj�]�~��D�qVH����~��E<��/��DZ�I>���V}�C1V��r�[J�B�b���c(��V��ym�wY��U���o��8wPO&���\-Nh�N�b�~5�o@�J�lY��{K'"	e�6��uB�����>s�FH~�%��+����!X6C�ɽ]�堷V�3oY��O"]�5�tE����k�/:"�p&����kt�`R|7'�[	�<c�p<��i�\ƥk��J7�g�K�����JO��,;,�CiHlV��ҝ��^����Gl���f����:f�]�Ŧ��2���j�����_z�94Xhٿ̓^����M}_�!�%�4��}D�,�R�v��o�=)�Lb!㢞�!�&����~���ܺ�-g��)� �/m�m=v9E4��	Ĵ��r�\��G��t-���Ȁhi��:G��Br����W�K[�E�5-H��� e��E������#z*�a��r�]
G㦪B?uj��;v�|A��u��v׶�s���5��"��S����[���"ۇ*��e���m��>�Ӭ$W%�2~ڿ����^6����_K0����f��T�{�f��aeuE��<r�Zp���͸���3qv��� �v�~5.�(����i�h3{U�u��νtl�D����E�&���^FD:#B���U��cE][��HlV�*���~�8}kxaP�ve:�`o\�M����!J\$e�mg�Fv�*k�]���R�)XŃ���L�[0���t�0������T�5�؜(<�MX�]�����Ñ^tA�s*�c�/B|�����ߔ<Q�)Nߖ2�<��P.�_L@`��|�!��Ք��*���}�$�-={hg�/�y���4�W/�6ḿ��G��� ������
����~�&�E)e@��"�_�ޝ��*���\��@��o;�	�s��	?�ຣ�\L�ME3	��$̫;R��/|S�͜��!��˘�Ve
Z�rH��v��ϗBx^�7ʍz����XRf˨3+�mtS�Q#T�dV���DX����C��:��A�$yM�29���C�^Z!�����E3˹��ț�?D�{~��������{��e���e������+/��� �fS�x�WvXO��tJt\_���k &�����tj����|���3�X��aQ2���`<��i�����򱖩��(�b����^])lތ/Y�Ґu����6WN�/��a�\��m�Zy���eb%w�˙~x�ɸnq�2��$���5G���p�?�?����œ��p:b��7Ch��]�e�[�T�Ŋr3��2�.D��=L�ڴ��
�'yq,��7��)<	��Cf4��H<A&v�%��p8CPiV$:��|x����Sj��1����9���KNH�`X���;��~ח�I0Znˁ���PA�f�)}�0oB5�~j�}����	X�y������yN��-/s��pK��
Ә2I|������ʯ���F�[�a�0�����j�Ҿ%\ͥp�u�) �<�k��������=��Ps���s�:7lŲ�n�s1�N�9#���4�w  $.�n}{�����3��&f�:x�B���3g� Glh�����R�+�xlsӞI���+n��,���M�>,�PL��۱�����
,�ҏ0��x�OA}"�U�Q�����Ȯ�۽a0ak�1c|�0r�w�����@m�]�|#��Y+�5���=M�L��? �п	T �}��D /��i�P�(P3�P�U�[�f�k'Ys YF�M�:���)N��:�:r>%����� }�%!������߲y3���x���e�MAFi&�3�K�Y�_�U����B����!I����I���fPB��(iќ��A���(I�>����56��Zh���B����_�?;)}�eƊ�Bu$�����䥴�-=Ȫ��⛗G�WI���lҏ9�`�I�L-2BO�����Q�d�4����K�ȉ���
�ꌚ��2 ����؞�f�V_Y�iğ��7��}��G�E���b�6��[9��1�8h��e�����[d
>xj<^`�5T���YW�h����Ȧ��r`�7p�-ȄFr��г���C���A�+�L�gJ��A��>�
�xlB+U����~OB�[�֨��d=���.��yӓD�lb�� ;<Y�Դ΅s���k�)�@�����Q.yӿ>�Uc��Б�Z�7�h�\����Y�u�S�}}6�Aj��E��ո%A͂5c|s��\�1��n_Gj�-�d�LS�2�}ޞ�\-�"%�W�������)m��
�*�y�W+w�`� 7�/n�P
���HTC+#���
%@p�l4�ݚ�=��Zg,��Xk��z?	A~Wq�S֎�^<ڿ4�P�*�hy�wZ_��S�5S��v��&�4W�|����)�P0�ܒ�P+t<�+��,HkfT��G�u��l�4:��h�K�A���X��w� m�jP�e5f��F\I4ZK�WA�Ɯ~����[��ȹӍ�$������g	�?�xhI�S��/}�����Bw�D=��"#k��z��M"a�Tc�ҟh믄>QV�N6&�h��|���#��%M�׷�CUw+X�������?��=*.�$�L��2e�U�Ә8#�e)�l�?�������|�G*Agb�6��3�ɴ�7:;���wؓ�wȴ��QH݅����/-�PC����l����SJ,���Vt��� t�~�B��A��Tz!�;�27�/�s��%�V��6Cf���rk���̟�"ĳ���x+
.uPf𱣺0������$ �/P97�}�]�y�G/^��gz5ʿ`���� z/S�.����Fa���oH�.7��ſ`��&�䨾n@�-н�@f�p.T�#oI9�g=�Ӎ�!����w�+g4�nعx1{��dS�I���=%�����x�q ��ʒ2C��%����J�ҷ�X��H�r�C���W�)��x���3�Vy��V��&� �,c�p�S�eb�emw~}fq����p�?�h++]�����HT���J�0}E6Ǹ�i翷 ��z�[���"+��um� K�nkȠ�il�	�!�5f#�~WU�(S�|����ΚX�,�F�Y6m���Ѱ�텽Ո*�,��%�뀰X	�7L�.?B�W�8����O�|J���?��D�,2|%�� ���@#i�m9��5CT�[�"H�����X�;�D�\ŏ�84v(�s'=.?�h�x�R�]W�
i6J��7U ?Ӣ���j�ɂ@� ��.PȲ������1�u��kv���߃��=�dѯ풖��Y��3����r�I������D�ʨTv�q�����A\spß <R� ��yg�
�o�r�R�yD���x./�H�lQd7��po��z:z5B�MpxD���V�Ld�L���a@ېw��R�#��J��P�����}0k�+�kn�9^�1��QLQIdt7�)�ܑ����*��D��b�#���h>����ֱj�b?�hՓ���8IV�Aj�{���n�ǍE��\�R3�N�gv@[?S;��O����RM0Ii���i�X��͡�Q�%�M�p[v���?�Ja��u>u��i��||��9 `I�e4��;�][\t(��i�n�D��t�8C�#��ߡ�#NY�Gf.�������I\�x�H��VC�5_䠁�c�&�3�����;`����(��&L�ЎHF��nt���rP���ͱr5�έ�	�������ݛ�^�?�9�1A���?4��1;�㴷65H)M���>�(At֑)��Ɂ ��`�]�x�$�0����R�Y��r�j���D�d�
�����6I��|��K��A�x&
M*���c�s�]�j� ε�<�+�����1�D2\l���Y��QE��+��X�ڿ�H����̋hC �2��O^.So%�A橂<- ɛ�30�n�]��*U��%!ҷ��a`�uA��4�����&\"��V=]bP���p(F,�/�~���Q�i���_���n�̛F*bET`R�I����=��j�i� l%�&�2�{��9	A��*ߟ,c���!y�|[~U�\�G.l��yD59�Ն�ց$��'����/�.E�O!Ҳy���[���ߋ��UzYQ�u(/�Z�9��ܚ0��ʦG~��\����Wa��9c��oJD�.�C��E4���>��'r%��n�V��	�9X�2 "����僫|�c>�z��+��1�Kǈ�{�مV"�!j���#�z���u�uI���Ljh_B�x96��I��B�m��M-�4Pj:�ģ攎��]��EQN�|&��l٩-�������Q�~�)��.������U�iB@�d�൧�'mXy)�>��d �|�A�r��Bb�ͽ�8_I�a�츖������P����%�x׺����%��a��Vo��*�VrT�}�	�i��
�E�]���0��*�L��vvH�&=���J�0��e�Vж��Ӡ=�X�5l����ST|@�w�r���ݻ��n͞+'�w���(���c3g`X#$���wZ�c�W�A��8�i�{��~�m�mI����f�����eSQ�grb�H�w�,�C?��F_���	#���e�sz}4��sfaX+ �އɯ�*0����%V��W�GG�~��>�Xp/6k�S�M������(Si������F%K�����
\i���Amm�&��l1kZ�;R�G���ʹ�=}�f<o�F9O ��ֶ�`�xBtxN���:��k���d�����zAia�M���ѝہ�:�f��f�b��~�����C�L<�݁��0ӟ�hY�Ui�4_�4�J}
�T�^��gS�X�������`�6�Ԙ���e��#�l�
îA����2� �N�,9��\I�.ϐ�g8���b��O���,릝��}�핰c��VT!�����1�S�dx�)1hf��u;e��x�8k ؞��Q��2)���D��k8�Y ��Һ��ߍ��%��Xq��	|�ꈫr+�z�mNQ�C˨��$�j=}]��K��7�ѯ�}�Th��ǯ߬�E�F��>d1X�[����s��y��A�Y0޵M"�{��nl�k�I-HK��Զn���8[z�<\� ��9'�Q�^���Ũ�-��d���½EAq�KH�K�-d�2�ZDz�����k71�@�ކV�'��53�����Z����b�>�ÐN�Glx�]��Uǁ�@Y��d��1T�<ɢ����":����5�M5V/����0�Êagԗ��I���s����	���w�{9m��T�2�KJJ�B��=��y�_t!T_f%��͸�=��#^��`=���+a�H��qSX����r0Kp�.A]SUڪ�f-�$ug�]~'�&��g遼�3{:6g���%̈́��"�;rr7N��ͭ
'Ip\��� m�h��7m�_��0���IgOI�gS�
�!��3!eH5(x�/FN�w�Ѱn�?mLu��ڽ�����_��g����VsMф`O�]N0WƊD�z�2��K}�-p_�Y ?tfΌ�##F��.�o3��Q�usx��ǋ�֓�Om3�o����t�?S�tV1rlQ�Y�2����b��NGx�<���S���b2C��\�M��@$'��Ϛ�tjL�-����C�"��g�P�~���G���`�MAV�!�EY���d�� ��7��T���XM$���	=�7�Y�,���(,Yݠ���&�9����m� ]Ŵ�h�'*�(p����g�+�k(��3B�#x�d�d~Y�?g09�0���!>qρ����M��k��ͳi��v��1��P� �`y�kִu�#V�v/*�@�(5/�,�E�l�p�X�*[��F�t$r��RLi<�#Ƥ;�Ye{+�Z��#A��H��%� y;h�G��fA!��_t�L����G�`����`b�@&o?ӷ6�͞A.����������Y�=f�x	���L������y��6��X���0�q�����S�r�i� �_،������#��]mU f$�jr�(��j5&E�;���G��&ɟ�C&�:��>���6����VF�J�p��:>�� �n�<�����ӷ�u���N�Y�Q�xZ(����Z���[Y�~�(P�^�����^\�=bv�xBH	";k�y#~|��G�w���K\\v>�C���|���בֿe�!;�[���:X
J���,)���F1���@ۤ+�i��_3�E@���R��b���s�~X~<�=s�NE�j>�}��4�(�_�|G`I�@b��pq��z+�k�!v�u�	�ڽ�JY�xy5rm|FC�UI76W��G��x�m�A��ӈ�����"��}��Z�M�I��.
s:�B(�x����j�=M���R���wzR8K�Tmj�zF�(�d6L��S;���M
<1X�t�I ���ب�GqP�hF/s\�xxz2�r���J@Y�\ȉ
�EK_�YR	�᮸�F��rҪ&������*�U��ڻ1f^�Z?��U摔�[�-���a"�~��%���Hh�����O^m�YzS��˲?�n����ôv�BH���3~�0��Q�(�����*V�</�tA��0Fŀ̔�F[�^�~�0�\�P�=���~�K���i]F~ة�p�(�3?XC_2[M����ɞ\�lˍ�E��� �M��>ܮ�z-��*~`�W� 1� �B���8��Q�P��Kx��0p��ltν�ĉW�'x$�������5oΩ+��&�~A��IUI�)�����J�RTʹs@��gɬg��tx��T���J�4�i���(���l�"F�3y�����(<`�˚<@g���z�ft�S$�0�!���IU�ܯ0�"��E8��%��4��Y]�ɗ�W�}nGZ(� ��_����ı��'��edV5z
U[��d��Jz��U�š���F|Ng���hʶ���^�G�gL���%��(�6A6���؆�m�͞x�I��[���r!R�(������EZ�,T�WeH@�Ew.����j��"ӾXs�l>1\����'��J��䵤(1��-��I���чO��mG�,2�tʵ���b/B�t2�O!'^���P�=��h�H��(����Ӣ�+����m���((����.PL�/�2�+#Ƴ's�B�b���v=F�Y9�ܾeJ\��X�@�e�#n�fT(RN{o�������]<�R�C1@u�!� µ�nO�]�~D*G�@(?;O�ɔ�M}�6�o��RP
�
�}f�< ���0�*�f�ZbK�3;b]F��5��������֯Y�fiF����e�H6'̎9,�%�D-��$N8��C��":�
��ĺ$=�-��4���� q*��]Cf[��zJ� ���ERq[��	��"��[�p�$��!��=�!����]O�xO�e�>��AE�+�RNH)����Q���=8�)�>������U��tg��[{��ɺ�$߰M��f��)�Z�!q�cb0��s���L�;�C����.��^a)��l*3�DS9��E|]w�zkI�)+#�Y��ےFj �m�}&��0�\�	JM�P/F���ap-�6;_�86���)0Ar�]s�ѣ" �]���\@�̑Nb�r�uxd�G�<F�:4�G&�H&GuG+?J�j��Un� � �e�R��]�/����1L�yࢀ����4T6� �oEl;Q΋мe<��Q��r�w/.��M��ϭU�a<�� '��i�2�#{r���搸�I5DJ8%:�{�+�CB�>1��at�2��^/�J
��
��=xB��r,�f�����E���Z��P?�c"#�N���4�=��u<`��y��>͢�w�s��K;�:��	ѩ�*�n)�"�U�s���[�����ӟS��JH��ͷ��yd�'2�r����1����&C�mȥ������_��)�0�a�΁z��چ�b��l5�3�n#d8� \��]O�"�� ̫߫x�/H	�33ԪWP���t}���^�\.���*3Մ-��r��5���"f ɰ6�!��u�\��p�7�e&������[q�9l����H]�����M6��Y��bjC����K���Pe4z3ت���	�V0^�W�զ5�ëOs�5�p�9l��.��h�6�I����7BQj���$���;T�.����j���y�@+J�T�Fg1�@J���3��7=PԳ`����:C���1Vډf�M���$,�K�?�	�����t3=�s����^3���v��&nM_�d��1���z�<��~�҃��񛅛DQƘ��V��VK��o��"嬆���sn)2��V���E��ó��f��#I�a5�nJ�	�U2��W�0�����y� �٢���w���;~���|O�����	}ի��Y��M$E,�PVCE*��B%R��� 5�a�n���@>�C������;f߀�¼�C��jl���i��tl�E������&�nAo7N�� ��V��N(��4O材��mv�?����Q�֊P�`���t5�C&��J�G���1˄2�L�O�Y΋gM���2�f��z�:WV���ʻ���v�ܡ�F� '*k�\�|�;ug��t�Ҧ�$�`�1+�'m۟�Ŵk�������˳&Ӄ���\�Zc�լ�h�o@���#�ُC����] tR
o4O���>��ޠw9A fK_d%�ֻ��������_:�7�p��͝�T�`|��=�W4�� �ѣHR��	��|���i�p�}X��yeLF�#y�(�ؒ�Hͽ֕k�� \�FA���F�KTN�P�JB���}J#[�툜�QT����(������,��2�;޻wZx���7s1	� �E�� �(X��<�F�A��+�cca��Z(_e���Y�
����~&d��!^:K�`y'����D[q�Is����IWp�p��{}x�q��T�Vh����� 靿�W�������u'�`� ��]����������j�G�V��l���ݛ��ڑ_��h\�)� ����e�[z��se%kR�a���U-+�u�	ࡵ�E��Y��X6���z�"�zn��1�RȨ�Y�-�kO��1������H�8 F^D�NX�R�k�it�ڌW���H�17أI�uxPQg(���O?�T�nbxA3Bxh��J���D�w�8��6�r��u���v f�FD>fi��5����/�R�����y�HR���A�������\��S�(�)M�"�lI�GȤ`R"}���ջ Lz{�8�ޮ$[����R�]�c��X�Ҵ�.��-#5,����L�Kf�wn�쓾-���Ǩ�g�-]�H"���8�K���
Q���CNG�M�	�z�Tҟ��yr������-�0�Y��*��%w��{�{*��,U?ʁ��fДkD��
�o��ҧ�ı�6z�t�e�uJ<*S�f� g�:�-�E:ߋ�&YFB/�=���i:���� ��g\���B�a"G]�PΎOe�����Ed@�ҙ��{���̃^T����k�
��^Z������;�}��$��nI�B�Ch�wu}��O���5X�>(IB[���QO��¸
�@����lt`$y;f8y-��)��&�	�F��?��&l����  ������i�8� �>|��Ɛ�����A�G����M���a��:�Xo����LUa� 5e�	�C"�mq��S����Y�N���ϲ""]��-�O����%.ύf�8)��eȯ����%��T�����q� �2�C2U�I#�[��*��I�ï������KL2�gԵ���`<��o5Z�E�xO5<S���֚&)u�|v�n�ݽ�����D�������곛vwL�&�n���JS��K?#d6�	
�h-�:=>B�l���ܚ:�bN�S�J�	�����	�>��\6ΰ���I렗���w���{��QyL����
�����F����8O{���h̴���Oӓ���/�]�-��v�E<d��"1�Tޣ>m�B���.���h�R�$��s���Z'5�"�֘q�Fyv�f1f���!�}GV�A��������]�9=��)�n��/�މ�!�#�1��¿]�������`.֕ݡ����?H�(J�����mjT�C�{�X1���}Wm\�_
<�A�@Ob�I����C��)����x���[��k^�+��Dv�m=�~TI@̝��J��#�D�vM�/���� o}�|���L�~����j^���:s}����&�;��r���!���������ހ� �ަI��}�MQ¥��q��FY� ��2�V|5�Oċx��=C�8N��I�`���&�z�(�{^�cՙ+S �c*�sL��xp�Pz ��Uo6�s�*�8~���c�� �皆��E~��l���8	�n���!=�$H�a?�ض��%�:31�� %t1 m#8FXw���훐�y�y��?7�`Ņ%���/�v�Bp	� �ܡ�"�v׻r�1��a ��f���nr:��E�Yf��:dܪ�^�;p�=2���ҴDP��M�#�A��+þ]#h��ȑ��i>	yg���ϊF<W��;�`�K���H�a�z0	��H�*y�h�� ;茧.�ʅ�aLh����g���bT<D{:�z� |���x45u��ָ�����n���S��/�P"ߛ �G�z���-ㄙ�P�]I6S2�e�1=)�O`m�зe@j&Yg�0\�ᱎ[𑣕d����r�./W�S=6�o0D��5���U䮥
���G���}�j1�@Z�2����:�=���1Z����jP=��2,�|10�!5	������Ruk��C�Nm3�,�p�R����M���f��3��J�G���1|Y�����Z-�ߟ\h�UV��_�V�۫�MŚ��4�O���|cN`(8zu$��͂Qe�ED���1B�>'҆�7��*hI~R�d�e{���7s����F
L{�n�yKcD� k��/��q/��ٹC��m=��"`�l�K��7ݻb5{Ԃvm�b�l�g��,q,�a+ߘ>P�`G9H���{������ ��8U�~����Y�G'p���p���6�����!�@�Գ��{D���arНԒ$#g�$��G-�����d�S�/(�?�)d?P��ʡn�kW�GZ�#5Q�"�ȟc$C9L����]<�z�"^%���o���M�a�
䖡��$��+s}^��B�X�a?�",C��%0�<�s�l��L�*���|���Q��b�
wsz���t���6�zA1k`�`���D�e5�l����W(�>;|a%����������Ƴ���k�J��p9��>1�/hp��z 9��Lp���W��B�@@=�/�����i�i
�x\"G�=v�u����G�ۏ\��q�r��r�6oS�n"���,��oB�`%{��mJ�Q6d��ҥ�b��a~!7ki�϶T� 
�#��97��q�{KP1]�����NA�@�$�쀖�S�ܷN��	�����SL(��wM�����uꘗ��\���/ !~�ے���/���O��op����A�ɢ��d�+������K�<�����-a��9w֤��T��L����Eg�_�M򩄙
����oPy��#&BM��˗���ޝ��.�T�w7j�v��uYu���S�8�:��I|��pW�.e���b(f��ӏ=�j�y��K�PL1̬�����痕%0�Kp�)$I���X�� �D��F�b��
�p�F�N5�y�)ˁ�����ȩ�i��P4T�;�K^�
yy��h%��q4��UOy^0,�=���ϵ#p���,��;@�Ԋ�̂�ܙ"�u-&v�[�)`׃1��#���z�
t�9��VN�r@,M�l�<�\>H�#_���FA��)�Z89 �� m��7��v��dDM���2?-5�����7y�S��m|�h%��ȳT�v�~�m/���/%�H8�K �\x�HO��u�T�˳�	�g�d4�l)S)y�|�	��z�v�i#fU����Ӂ���n���ƽ�0��Sl�A$���b�~EV0�|`��ېq����'���׈,�A�~��NA"���PLf&�dl{*��4$A��wA���&W����`e�VC��*5$�%��,�6��0�;#ʀr�� ��11��ԭ[��\~�}*�IU$�U~����:�s��薀�dRl,�
��w��o\!;�tX����7��-\�:i��a��& 1I����Yd�knV���V0qx6mٳ���ޚ�_e;ܘD�C�y�_��̮��q�p��!�S���cQ��&E�Y�y�<���Ǩ�-��?�9�`��`Mި�&�f�A� ������G+�AEfzV��ܹ*� ݊Fʭr�'/$��F��c���aP�J��I�����u .@��[j*�Ab\�r~^HƖN4
O���jK�(����F�yގ��'UxRB`�G���]�`��(֝m�inkm�.l����!`��:��O��0^����hx��>C�
�G%��vkZK�k��tQ��w�l�	�#�Y�X�(��~W��dy�@��`W�I.�FA%&�v Y�D�]%��݋�R�B@N�P�R���WӠ�a�=!E�5�*�d�R��+ܹw�9^�F���r��WU���p�{�����_� ���i>�����j<5 q������_�'}O������Ǧ��^�>�$0c�n��EPJ���X���FՌD��^��V�@2g9a
���!聀�B�
�P��'��IAb���>�XB��T�Onn�⥋G��d ��9�K�k�D`�D˲���!�eE�/ў�b	�t��N�&gU(>k$�$�ҟ�{���Jm�0<�:���E�҄
�}6a��.�er�}˩���t�2`Uֽ=���P�c�)XG�=.�6�/�vua̯ɘb�Gk*"��i���%�� �} ����&��BE��dR�M�4��>���:z����N`��t ~Y�!櫾#B�H�_�R�(9A�A����|傚W�����io�&X� ��K����W"���g�Ф�[�����=��I����JM������;�|�0q����e�I��!��A��i�胎��5�z��6p�*�ʔD���q\lÀ�ʇ���D�d��7d���$w��u�J{��D�mr����}��L.�5��*t_ �w�#��E������Y�/~Y5,�S*B'����z�$����W�j.�i����U�s*C9~�J���ݿXﰥ���4�~���z��N�m�����Xr#b�\=�����$5����j����R�zx�裏��#��U��|�`^����9�*aP������C���)\����d=�_�I��g8o�튲�O�<OD�^����B N!�ľ�듽lX��N݃�T:9�~K���j�T ����9'M���WH$xD��8Eb���0���R�
wbz4p9[�����:�a+�Hr���� k4I�<��{� "�zF����I�(����kR�q��m�	�u��	��ѭ*�p�	*����4[[�6Q�!M�NC8tU&ǚv����(��Z��Duts뺯@�z��.1le�fH�w"\//f�3��i��!	���i�P�,P�gI�9o��v'�-x�6vл�6�I/���27܅Ț��_o�j>�cIކ4�è�hϜ�-�9�t�}���S/�꠻œ,\���=�rb�jB��>�O�!��t��w��AO�c��ݷ��r���O����!����2�F�|56PW>�%I o�_������o��>��!:����ʿ�&�^�#5yeGf��OE�Po6���J��0�y�^� =�Sl�ZSh�ӟp�[�f��f��{�EJ���k�������#{>y.4��<��+��g��Y�^� ��ocj��2��5�uZ`��dH.uO48�~ T�ŗ�e��\:z`�+��)L=��ܳU2Ol�5�X�na瀤�Q��j���Q1����X&σΝ�d26�}djC} q� <�.Q{G`t�ڒ��0y�Ć[o��_(d2ƫ�}	5�I���1�{�I)�sH9?Oi��K_���ٴ�E�J@N-�t,HD�Z��r\�"��0o-4���(
w3z�%�kP��Qd�ku��ܜ{X�^��1�A����Y&<�}|��U��6�děr��SSXK��+H�@�{�d�p�,����,���`t�y'��L{��s��g��&sp�|W6p���VH���ky����>Hӓ���x�.��H#8�TP2��ۯ�,߃��f�R���s����u0��(-��2��#t�RQQ �C�|7�dz�t� �IǯM�+�����r4��:p�,���+OVmb�$#�޺�o�CH;`W34�ob�%���;1��_��M";l�gQ�6�ۃ��p�e�x63�t��8��I��Z�?05��:�,���pAsZ_!l�Jƭ�v�l��纔1$� ���9�a�0�C@O-X�	J\�VrCòuju�����J�����U�w��2��W.!�q��.�DJ�Q��S��6�P���W=W���y��W����2N˪r� '�>�HdR�O��^b��N�'��f�@����.�r:NI-�"Ρ�U�y�#�Q$���ao�D���ҧF|��T����-,F;��/l�]&)�w���.�kzD�P�&X��9�6X*�vo�����<�A"����?���p���@h!˛͎��E�1#���W81�!�tNb�y㎞h7�Z��$�u8�k����Xg��%�����B:�8ݠ�ؚ1�����NX���ؑ-��&ξ�'�{-��
���03X������Ăslo��0��K���<�3`����d��ڴ6}4A��Q���Q�bQF ���}�/� C`��
f:A|S�����i)1�]�=U�� 
mKam�����i�q�����lz���������6^��Ss��M�#uL���e�N����x,s�U���JT< z�/�y�Յh�#'T��S�8����3��T���m�� O}@�t�`7��ý%O<�)��ߠd�P%ȟ���"IlN�X�a�2����)B<�����%�N, k:T7Έlނ�V`Ё��]��6�1�z� �0AzF<6�8E��]st��i�_��:�_.#
B��}�}F'<��DQ�� ��%�Xaw�ʬ)�+��Am7}s:V5���ΧI��������ܶƗ�����m������5�>`���"h�X'�|�6�k	�asIe-(�o{b.o`m8�HT1.�{'-�0.�3�!ӭ9���:>h�j搎�Erk6G�ݨ�|�9�~*h�l�b�*��:����_b�e=`仒�gP��,c�]�XG8�4�z2�ŗ���*�=�-U��]��Lq&+�_��(����m���K�΅X�Ю99����K�)D'�dJbMd �7T�����q\��6���m�9\���`/|ў�6Y�U�h��鷜 ����+ I��[_G��O�������վ.�D� ����ck_�HT#?Rz
2�%�bm��E�Q�z:�7������x��c�����g�����ةB<𢨠��о1Q�m���sg�b)��°�����fL�e���ad ��8n�:�s��oy�z��f� ��)R�f��S��R��4���7���o�vu.��߶c&�%�.xL[%��?
�Mӷ�1yD�и��Oi��;�__I���8؀�ˇ}�~�Ol���W�)c,��6AE7�Q0�����jfÃ΂��Jr�t۽]m.� ����߸c�ɿ`-��\��c���Gu���q΋�y���A7���?�Ѳ=X��ԴtW�e-�����9�W��f9�0����$��'�>��J�d<�)v;�a#P||P�!?�j:�C3�h"�^�&ڜ�SE��R���+@e��*��h~�/��gf��$c�ߞ��8�0��&k�!<*G9�-�M��FՋa��jRK�Sml������ ��[7T��rWn�l�О����+i��V�E
����٬�G*y��2�����wͪzrf�/g
��7ǋB�Vd��]�bx��63PQ��TP�&�]��k�e��z����w��/WK�7.�[W�d$�o΂p�)2��H���F<`�*��Y��c�HԼ
Z��������_<�Z�3(Z�$a��<�n�wp��k{�z��~1ZW��]��n��q]K��kz��j���HU����Ӭ'����gb����l�z�9'�e����?R��ZlH��p�\k�]�1w�٭���������>���0\�@�6n+а�č0Ly�T4��*�(������r��ڏ\��(/�4�u���!>���/�u�ޥB��)�W5�`Y���3���d��V���j�VH��ْ^=��Eg_��]G��@h�;�̾l��m-�O�T�SW��[_d�(�+���޲��f�|�����HW��N�0�jm�B�����(��}�IJ��^p�:"ٝ �>���q���=�d��.I�̟yV�k,�}���&;�\6H�xz_�Ojٙ+��jqr���з�T�р���7�Y[%�b�$s%2�8��3n&u���O�����k��:����'�<w�o)��(��m
�9w��c	�|�N�d_��O���Y��60�Ш"mr���ڳ�{$���0��V��?n�>u!+ᚏS����䇖k�k%�F������J�V�+6��3�Z�Ո�i���P~�M��ǌ
�0��r���B6	�w�G�/��k�7�
YJ�i����!I*�m4�F�Ţ��'nj#�5�I*�U�35�yӜ2���~�:�9
P<�m�jb��J[�i|y�P��?�[�@e�ӏ�1�fw$�PHO�nks���3B�ăc�Qx�Eޤ�X��B���j׷�rNrEiT��2I���E�2t����8gzm׍��fǷY,CB��ز�%w��(E>��� ���>�j�"q��FO��]�}��V��9]���{��o��O�<��}Jw���3vlQ�ꛊ���Ը�U�ھ�OE��ɨ[l~sݴ��͔�{������v�������Iƻ4��J)�.#!�(�W��v��~��Z�ȗA&��e}!�����>?��6G*QH$�W��\�����Suy?c}w&���k߻����l�`j ��]�%�\煴ƘOh��=;��-�5���W0i���S�ɉL[�ԺU�Ȟ-�	��Df�$���:d����Ο��h����U�<������w骾!^P��d8��t��� �*W����l�b�"�sda��;�xֹ1 ��^㚅V�Nd}R5�Fm"��z�p7�( ���
�� ��A_Xh��L�`h�x������dJ`9��/**|ʚ*]j�²��S�y%� S��Ҵ���S��;�=C�q�
rv$.���7k�A+�^ӊ�A S�u�_c�:@�o�M6���NT�N�J�l`װ{�sɠ���6D�B�o&�3����ƲPh��ʹ��	���V]�`ٕ4c{��.,`LQ����4	����pi��J&�S��3v�ԪA0w��zaV$p���u�)���[53�F���M��4�*����O�و�b ����G��q��<P��A���:����{]Z]�L��x�wƞ�|(1��/'�G�XF�(Y�y~���%�0�Tp=��M6��s:@���m1;�P<��*�c�&�M04ztΜ���]S6�<9���|�K�#�#�����	�Y��h���m����]3�[rf	�y��ł�\$�K��2)�;,�}v�Я"��όq��&�%c�]������q�����b����%�t��˱R��м��� ���F3�L�@��� �	��O���/�P��uj�P-� B���_dK�>�2�tj���3�1W�.�%��[ H�ݓ���{�f��5Y���[�_r�r���?i;�JY����.L� >�8��ߖ]���K'�R�� J���|�%����9v�O�58H[?�3�y�ȁvsT�I�G0-���p�{Jn����h�+&��E������F;�h	TT����&N�Y�ƕ"�����B[��{� �+ӟ�k��	�H)������ةGg�3�*9 =k��?<�୉��>��8F����Ii$.���Ա��_W46fgI�����\�I�����Y�ib��m(�:��{K���ύ�p~&D\��DXg8�2�G��k��[�����t�W$DһIF�7̰�bM(���Uch4�C��2+e#�CӘѲ{�h,k`:�F���iȺ��5�s�Ζ*�ϰ�y�Z
��3�8�^c5l;W�vv�	T���SZV�]��e���￪zϹ@�_����� �2����'��:��,����E�;��榽����G[�Zׅ	�g3��^��w���e|j2� m����hxt�w����Q]���v�S���Ht)���Kv��	fҧ%/]g���uR{��mEMR<� �Ѥ(�A���*́Y�ò�U�/(��ь[�J4���r��_f�/��N���i!<{M�R��Nw�(w+r�6%�X�$�U�W��H�l�/��e	R�0Qc�ͷ��=փ�ű��⿦{�t/<�5��i<��J�.*8UKٝ�����w�$g�ԛ�����S���hmB�]M%7�V�F^G#V��m�2���س�lT�?�\�����)՝�J ���>��[8*`X�-	 ����5��c�.��f���L�l �\��	�F襖���%�p��@�`��˟�{���Ic�=:E��	s�G7�2S��1t�f���|V:&5}i�EV(g5[�^2/�`\h ,!7��o���V@�(�{9R�ċ���^,�9>7m��Ӯk��	�P�bK��LR�	J�g	�&\Q1��,D8Z^_�����`2�"�W_��`s��D��+�\;�1{*��@��T�S���Tb�P��������|5�.9�3�a�é;�]m��T���HS�:��S܃�XZO����0K��z��2rc��^�p����� +?�ў�O�ω�lw��nU�(��p�Y��+��Y�R- be��[�Ŋ��G���Nқ�x�F��o��� ��¢��NN�E(a>���u��O@��%�9��V�1;�k��S���ԅe�B)���I�X̹�*��M�����{ޑ!s�#���(�-��x��
lVfHq� 3��oѫ>�ߡ�K�كF$�M�1�cI�S�K�y,��y}��:�s{Q��%\�L��K��{�_.�h�e� P���@[�XV-=ި]�ԿT�Pg���֘?t�Ś���m���]��,G+،������fc�x�鵮��B���l�W�3�J>m�w�q�õ�bp���r0Ts��AFLr�;9$��������s}r��f�<X����N�ϴNV�PW��<���4ׄ��=Ah��9�!��3�ŦBGL$,;������/~��*+��"�!����G��X{�}�x-w�z���c���-�%�{��dީ�<�мQ��_5k;׉xG-���z�u���x]p�-���{q[[��l����k�D_�MA���_�����|�!�c�+�D��8A��!����p��M��0���^j��i�R;k�X.r���hM�/�L./^$[�1ţʟ��s՚fM���qVH8��0�K��1���i�S�h5�����2����RVVRᙑs74mr�X6B�۶��C�J拓G��c�,��{��}'�4&�cA��\�n�Ɲ\�e\f��!�&���s�u�F	t�$��Ϯ�O����p p�@�y��HT�ҩA=����В8�䷹�țX��񛕻1�0����h+s�)�j�> ]7�S�`/Ea~����M9)�����ȍn���Ǽ���"��q5��yE%S�6��w��Gh���N��|pC�BVs�n}P� "��ԂOu�p3���ˀ}�\=�G:qF�P��t�b�.7�P�wjp&����F����>9pA
���/
[eJ��z��X�#=�&�m���i64��L���u��}`,3:�;G���Fr�S���ik��B���Z�|+I(�IJ�U~R�b1!�C[��P9 �h(��($8�ym%l毡�`3ր��@��`yH�7��4���.����M���\�f���Ү�aF�t���f���ۘ�'q QE�/_�&�kH������xF~��D3 !����.������qJ9��Ο��ذ��3��oe�W�h�^[�����P�j��tHX�H���%��ϖZ5?�t v�${, ]�lD��yj�<�Q�	-�H��n�x9&s$�� s�t�����j7(�_�Sw�*�ӭ�M:z�]D��T\s`�8�{%¸�bG`�ι��Yr*eL������j���z���!��3Q�V���ş�Q���V���\j��NUV�2�v�q7���5�)���~'���5��$?yG�qgV{��\���!�>�mv�:�$h ���B[����#zoܪ�chG���o9JK��1z�-�[+/�٣���b��-��=��c�� �~Y8�=P?��S
;%do|�Qt�0��Uכ7YO���T����	�"�@)JB�b��$
?z4��c  }1�93�S��S���
�`N	���K�-n1fܜ��)xDv�oHv)Z��%���c��{���>-NT\�<j��;����R�2۽�V��t��r��7��P�Hu�/�ل��}�#�B� J�e��X��i�Ԉ���Zt�4����ݻ���K2�LUh*��<���;�۾l������Ia��;U߯S��Q��3~d"���/����7T��Gy�7�7IFn"����*G�Y�tw�Z��3޸�&{)�<��;w����"�5���T�&'����^�zg��A�ȽHݴrL"�Կ�Q�Lf�`��ߦS�(���M�3.��"�d]�����9@���p_���W��JN�F�N�-�)���`���l��l̩U�{�Q<����G�?��s������u`�L�yifC�������b���.�����!/6���0���?,��n4Se�`!�C�}T��r��v>)oB�Ek��m�=��%ޠ��2S�D��0'kA>_�eHQ=��HF־O�������^������V H���q�զ;�J����`s��|P��a
5 (� Ʃ��*�F-Q�@�{��<����NA�ӻ1�JX2�
��t#>iVxs�kn�!1�݂�eX����ZB�"��J^\)A�GX�3E����c�/p���n!Ь����O0�/��>b
��Z���\�?����Õa��js��{��>��\MTB_1�5(�(VY)�WU�O��Lc%�ψqЮ�Σ�n���Q):W��6��Wx�q0ۃ����?�����gE�#�&b�_��*)�7«	�BZS}����u�b�l���Ų��tz����j������%Q^�9rEl�����ȩ�w q!�XE�kq�ɫq�����8y��S� $e��}	+�~�LW#�A �5L`�W٩}*�< �܇��)n@��:eg'e�D������9�,}����A�;j�s�⇥#m�Q�I�����-���e�2���CN`T�ߟ�XI�}ZY�2)��1IH��mYRe�����;w@A�I)��>*"�c����&��H�����\+Q��>���Hד�I�A#��BV�4��D,�4�}F�O��78yuj�_2�=7@7��.^<{����!{�n'��/i�ZE�w�S�LХd��pQ8�f�/I������_�P)ǭ�/���f�t/p(k�k��@���j Uf�m��}R�^�+����Ј�����ós�<ǔ6Ԟ���o��>��h���P\#ˉo� �Y�w���ڻ��px�P�:���[qԝ�Bzv����ㄸ��&W��_΄�͌����>p~m
��fS��D�Z������uT�|p憽�F�n�����d����0�Q�Ņa"l>1����`)��F��M��?�є!��L�/vv���,�W}~�����s��P��w�o�9����� Y"�9ȥшĿB8��(GI�el2PXn�mW���\�R�"����Kic��oĆ�4��HD�������+��ԓ�sΤ��::�=�[8䟸J�����F�n�+T?�]H4wҤ5=�:����m�C�[�����X�/�A!s�(�f2mw]*"� �w#%n��n+����^YS��rj���>u��۠r^F�z4Q
�m��8=]����'t�q�i�ذ��s�LS�cy9{�:�H`�=>Jq��i9���:d����Y"r)����T�>�~Ku�[�}��=�i[�^IU�/�u���R�n�)`mt���g+��,D'��xuwߣ�:o}g
�� we��i�߄�ĮJZ�c�H���|XV��`��
ޒ�*� %�Q5z����أv��!#�u$ H2���`2/�̬8|E���}`N��q��Ԑ�C��b~M��*�ƈG��j�� ���'J-)	Ή�%G� ؗO0�0{M��y6 ='c��d�����Ai��UJ�ZVxk��$ �C�0sZP��g>>)Rx�"}�ި��^��LnpK��8�����:H�kQ���eS���r]�;�+�PP2���p�o鮸cc�q�Ɉ7�f�.����@�{oa�G�= &�2"�&�a�+��AEI���2
 H�&�x���HZ������	}�m�W�y�x�Le����Ou�܂	�}3����u�獥V7�~��Na�J�@�;�3��q�܂l2����n�-��e�˖�P��huG�;F��%��L�`��);e$CV�Ԛ
�~���4Y���Cy�ύ�E^�]|FT��郥�%:�?��q�=��TϮ�8���n/�H`���Ȱ� R1%ԏ����z�"�� >T�zha%G�zzu*H�{�3�	�sU?Š�lj�_�%�Y����Ǥd�_,/ <;���+ZG=Y-�4�Յ��o;�B�!�V	�}| ����*�юk�SD�+�V0�W%hT�0�\K��+�#�$rϙj�Z�n��ȋ:���.���(x�/[���?I�-Zܤ���WS���~4���,S���A�bX�P%��?m�6s���EN
^E7+���� ��3v�e}/[��mC�aY�@� 3m}����&h�ոر]���ُ�MrS�ޖ�����T~)$�+ሻ�G�7��|������㿇�`���I
�@hW����`U��CԊ�3:����N�4<��<F݇�͟9,3�6�US�h��|��H#%mO���2��R�9C9���#�=}��G��m�R��䀢>�N{��k�����`QkV���m�f��F�{��:�&�;�@�F@�\�uS�|%��},��)V`���7�긂�˹�� ���O-��q.�#��`!±�.��j��75��b)]�f���d=��4M\܁��c���3���qT�&*��� ��|/T����=�xB����{3+��?8ǯY�婐I轺ȣ�]5K�嫩?�Q�c5w^�j%e�����3�⌥G7���^�j���ޕ�z�~eǸUq���<�����Rٜ��-��yyO�M=������1mu�l��ߘ�R�Tlq~�K$*�!���r�뺬&:M7D�lt�v6X�M�
�{cҁ�l��"O��,Ze'���!�@�ݎ��{�J����x��v���#�k��tJXT�|!y�����3rx���1�[���( ��=��_���]	�8 Fq�����q�>���;cg#�6��3u+������H=�T3�}
_{��N�9i�`�j|���cB�q��8����BCul7X�L5�p[��FpmU!�TZ1�%����u���㮙Yo��R�?�,1aBϞ ��B��`������h^~�g�yY	���8���ֺ�� Gm=MJ��:�>�cA~��?10Ql(���<_I���,ZR���64*�b�5H��ݐ�ǋu�.�d&�����@_�����Xi{���>.�e�:U�˦q-o�d���zƨ�m���G�8�Ꮝ#m�*�(F��pq���0U��Z�V�gI�1nzĖ�lg}#��V�����hf=!5p����00�e�mմ��[f\֗ ���Χ���]���a�`�S�K-��)*��>��v"C���0�8M�Ju45&�Uk��S�m�U��Ρ�77x5i���uFٿ��ZsE��h���n����t4/����^��׉�:��?y0/��tN�P�vh�q/�AdDQ01��3���[X����@P����v720%�.R��ڡٖq6�z�h�y�K�BY�ȴ����}:%T���bm:������`g$�}3 x�f{h��״�cO$�!��7���pvv��e	`W��*ѸK����Jnj3>���a] b`Zj��?�UՁ�e~r0�+/n�J"���Ψ�1Oa��[v�EwD�d�(��z��5���T�V@���4�bH�=iZ��&bh^`l<c���)����������q+Uc�(�t�� ,�
���1'�͎n�)x/���L9� �i���Be��n@�1��p��{�=�ָkW�ҁ�ٴD�0��|P(�������$ps��PHN�$����D�k�4"#6i�����}�܍�����6	�8j�1v8�@�次u)�2 仫����/c˦��F�|��rc������R9,K�S�o+���tw5f�I��j�s�`3|�w�3=fr
#�Rd���4Z�f;�X#o��B����輠�G��"QSћ���aջK�)���
�G��S�,�;�B�f���;�.W�>�\Q,�짫߬��Ǵ��Q�'=�� w&��Ԟ]����!����+�	�Ҥ5�i��j҇�U�����<��{0�G�������V���r���R�ɏv��9���UN\M��R�?��Ȗg��3d������簿�R����J�^_{�I�'���� �S���]>ݓ5
��MW�ܕQLI�(t���:ǖ��m�>��<|Z������?@���%����I"7i�Pv�5����x�$x�_��(��?RR�] �9�c�d*l�1��'��B��W�����a�ǎ�&�m�7n�B
G,�_�ˆn�.�O�k���ɀ�Q�c���c���!�H�lGpli�u[��1p�@�*^�����������!ż��z��"�i'�p�rD^}�e���hE~뮋����S��8�%�zw@.�ޖ��~�; ��b.N^?Q�*P6���Z\���c��RN7ٴ_�@�ק������ӱ�cͅ}
\��bnP*\ͨ,���pR +VC؍��P����Qf�;�/�vp>t�\�B���P�ɹ�i#n��L
�G��/'�l/P%� �_aɱ�:�Fx����/�E���*��.k�'?��wG�$Uː}F�K��W���?�2�r�:V
}�k�,vL0�A�A�qPrM��p�v�>�]���i�P��8�� �_�i��{5�Nz䁵���xZ�0Ė��cw;�F!$��F�6m8����4o�@38�g����*#�_�bw�8��H��Yڢ��6n������@Ϣ�%K��t��K�<C��(7e��Gɤ�@�'6��{�BvMׂ7��� �,����8�3�1��E"1�rG��!m�caM9ҴV{�̞�C�ew1�.����*���oGo���H�%A��k<0Q�;��~��[lމ37���Q8��NU����0"��%�eKJv�sˬF"��u�M��^M�L����eU�v�@]h�ۧ��~�z���~q2����N����%���t�k
AJ)F�#��aǝ��O3�;5�K��u5X��"��J�[8KWm�?)�?�f�����g%�M�`�$*R�y��=�̢KNJ��&��R�5���W�M/_{΅QD��	�+�]����Ь��$KLgS���U��bd[a�����h����f�`��VƠt�=���<�y�w���x��0z@9@� Wx4���K�/~I�f�Wf{������'T@�t�x�YV�m=ؠD@t]&����=ۋ��+���h5Rgԙ�SK�=�Q��2�b�@��B���kt2��4dU~i�)��	@�!=�Es�����;��]�؆�W�����^�S�.ub_�^��� ���t�=��p�rz�\};��� �&~)\�����ڶR:Eu)nNZO�y%!~QO�	��6�Ҽ=b��W��b��r$�q���ɣ/���:w>���L�Ơ�=?����B�:�A��9�.��5�]�]��ҫ�)�,L`yĂ�$�xڞ���B|��oO��������G��ܬ��$��&�Oȵ�c�1�Q�|�}�u�[+��An���.i��&Q��c���M#Yb��a �˜���H�e���֗�CO�uJ:�4d|��<M���Vг_�/dU�O�n��֔_�­���(���l��[�>*X���a ���Y W2:&��p�Ȭ����v���`�A���A��i�O� �����
�A���o��M��iw;�0n�6�X\/4�����=a�$�r��\�� �g�wGͅ��Jw@��O��ϫ����o�a�%��|N�+��U�|��a>���ZP��5!�0k�J�u6 �(�Oǔ���bvR��O��n�J�5�� ���������oY�#"�XCXŗ&)��qgaE��c��WvQj�X�BJ�SGS`�f���F��@&b����9Pp���q���:� �L�g��h�%9��om`�����f��\�.�H.����s.�?��<�H]@-���܏c��L8 ��6䋓-GN|"���g��Pn��%��ړ���# �A'ʀy�T��*1�t 5���a+�������M
�?GuCU��Λ��=���f��Jv��������jTZ�O��B8�b�ϑU}���z�>����m_���Rxil��U�_K��ڠY-�s"B��$�lxߤjsx��.8y�S��j���@ɻ�V��+B��d����\��O��F"4���<�9��ln�G��#tx��q���#��$	c2Y-�UH�ܶ2�U���M\�H,W��4Yѫ; �A�=�D���lY����F��o�N��uwE�V�%L�^�"\0�^,y�WiD���x��G��������_K[�!a����=ɭ�t���� �vb�N1��F;���t���蹜}�ߓ���`Md��\���K�'<X�VBފ)QǸCm �h�ǑGE0�ۇl�u�9�eiy�h���Vc{�fn���sU/���u�9���(¤��>�&D^<�}�7c�^�N����/�#j{�}3�6��n�U�}T�Y��)l�'��"�#c�(u�3S4t>2�I�2��/ϰ����R�@�V��� �@&��6�g��10"�mج#���gC۫Ó���RPM�s��#)}2��{��E�g��� ��LQ�`7��Zȹ 
L�R���$)rNo�����Gx�8����0]E?��p�C��Ċ�@�ml�\��CH��<z�'c�%#2�ٴy�4t@~�<�(f!I�O!�r�c���-[�W�7!��D�X�uhV+�^2y*n�h�`>|��y-L@���0vڙ �>����{5��ų��w|�Q ���m�%�K���E��*�C�w�(�E,��MQ����U�2%��g��69z�4�#��Ԭt������C`���AD)֕�-����^���2'��?-�>*�ӧ��ǝIA����O��Fγ!���!:�J��Z}d���uC0�+����b
�)Ȑ7c����쒍��i�:�O��$fS�/���_��@�� �<C�:������\���>������C�(��d�s�BR�/Uk�Y�ƚx��/H����Ɂ�҈�ZG{�����休4��R�>�&pF^K���V�u3Se2l��e&�*z���΁_*�ay{�i�X��;�L.�$a�YIWRR�"
�N��%m�2��=.z;mfSg�>�Y�V��<�3`^�L�7�j�x��p�n�Ē^���XRG�ˎd���ܛ�������:�X#��D�U2�"��?Thq�GsZ�=䭪�r���y��O/��L�p8u�@���sD�]�T�HV�LB�9s3 <\�����O��	�)�R��Pv��fۡ��jPާ��#��K ���3��w�1c5=C.�����jxŝ�(%�g
�B�ز�
t'O
�êc�����B���x=�)�'�d��,c���:��2;�����G=>� ?�L�=ؕ�t:%"�P'	(��M�'���^	��+��/�����KI��u�K�"��Q#��(5 �WyS>\[_�[�U˗8���E�/����B<*��@!�F���{�{��ů�:�H@/�~	�0[0�3P{��F6_�������H��kT��$1�n_#���������38#�@1���T!�%�� W���m�}��0D�Y��ЈnQ2z2|�hT3��j[�4�#f���j�3-r�Hb�)�P��%�u���h�N�Py\�X�,xB.6��-��a�Ĝ��N[Y�)�/�I�%���H�L��h�ǰ��v�|7/����	Ҟg��1M^_����Rs#hO���Ǽ̦���M�Y)�B�Ѿ�lO������o�̏--����yz��ݖTyH>}�
OD�=��t3z��#e ��l8`%��g�|�T�gD�[l3�i��NL'j����)�Ǖ"��6��`/�/��*�Vl<p��b��'�D��NM�>Ʉ�۴b��\�fJ�Zj���l ����[�ɰ���+�\H���$���cyVp����3q�����gJ���Tɽ��xJ�f�3O��j��HHth������0[��:�zZ)0�ukC��c���Y+�U����%�G�(@ �c�0~'���6��S�+����X:ݿ��H�}�Cc�w�	�W.��TU֖��%����cAN��,Ŷ�0�u�\Ƕ���]�������C�hy��k!k~������k�����{��$_Ț��&F�]w��z�T�)�Ũ���D�e[�����s���{̶��s_���s6R �@���/�P�q�;��Djq�����PL�R��K�7�������9�nf��9�4���j�+h3i1�u[A �-�25^�Ym:͢�E���-٦�y��s�ऊ.�*���g��D�#�^(�	A�?O�K4��VX�T��-`X�.S	&�5d�-L4�Äz܍=�������Z���[)���}]�n��k��!��`bpn�x �؆��n�	d[��H����<�_-����̌I����1lC�ݳ�!�4�&Z��KܩwVs�-�ub�s�I̜�.K���L��ʲ�����f�x!�M�ۈz�? 2��FWh2�P����I�#��b��j�|���E�A�HO�lK��UA�R�e�>`ݤ%���Q���V[������a$�������%֏�6���E���|-ӾTE�ÅO����o0{)���������w~��
�%��Jp�ҠBd�l�d�����jWF=�p	�v>R��H�o��/�X�!��Dp�<�ګ����k�p%+�B/~d��-��<wYr�EY��q���'�c,�i��b�ī�E��C�*6xml�;�6l�:@�X}�p���{�<:��70�+r�>X��ȆXe:q%!��΃��p	9�������.�����("��,)�n9rG#�����W��nx���A�T�RQ�T����s^7��x�o��s��%'�vM��vu��0��׿S3�a��R�֞K!Vǒ�&�2��Y�d܈K���,<5r!����=�����l��ϴ��s��aJq(����II��{����9WK�X'M]��@]	~h�Ӧ����F���E�h�s�O�o�h���S�(�.��v7��@m�R��l'{�`L����\3G��3X�ٳ쏽c��!?䅾�و+�9{V![K�L�����Ĳ�n�dן3;����6��h;~ո�,nq��$\V�`��f��(ı紘�L���������*[��sP�S�ܰ��j�"z�8k|�o�M� )�)i�g�=T��[^k��7Y�(�u�ٵ&T<ʹL0g�+T��n7U�H�C�a-�C�,�~7�� �#-�d����{���b���c>�\�P�L|���U�J��Ą��u�* �0����Y[%������u�c��S�}C�X�����Ju$?Zgfd�n�r�����5�;���:����!ۂ
͋�m<�L��6�;�?y{���3,i��WE�Вz���v�f�r��f�p%�� K�C{KA-+jsUPՌLP�%7���X?Ⱦtz�3��'z��$u�gg��EwE�w�-���R�8�n�/��(p���+Lc�[����6F�S��u�g+(���n�Bѱ�{�{Ɍ�Q�n��	��B�u��y_gx>��Қi�Y���N���I�uM���ct#(X���n���Γס0ʣ?�"��s5M�K?�6��]�����+���\�mk��ִʰB���pN�j0�<K��#آsK�l=�0�G!Z
��ݟJ<ݩ����G�1��=G�5G3��GU�[��x�#�0�۬�o����~�x�f�C9W���)���@)���@�@��������-.3�.DAB�t�) ��(����v�{���y�LU!~Nl�����N|��S��d4�Gc��!g]�S߅h�4ڻ�q���1�0�S羴 ��ZٸߠGsHr��.M,~=�m�48�i"K��l�S2�z�o��/�l�J�1�|?��V�Y�ۏ�߼^��'�pL�Գ#���eQ�v���Ԡ���~_>�#�� ��Jf"��̒b�����+�5n�A����+!�E^1N[9F�ܽ�e���(1˫���.��5�$Ǉ�o���-�)���H�.��T���[e��=B�H��4́t�
�5ĸzD��c]���t��|�Lu�o����]�QHo��d4i T�.��r�j����r&�������:�C	�X���'�U_��o��j@e�m�)��4d2Z[/���BJgx̞7�D���F������H�9�,jq���6�ǖ,,�5
.7���_��8c�p~����[�̘������ 4ks��\��
�ot�<%U% ҄0�����_O����>�S< ����/3��^�ƷBD�n�\����L6�4�@-�[k?��`>S ���?f.�|>ǅ#����-(~��7����v�xal�B7�^��3�<؋�����XbW5`.%g~lq���2�cYu��b�:�Y�Tn=��^�~Y�Ê?�AS�����b��`���i��y�P������A��$䛞�,Q��<��o}e�Ʒ�i<4���| F'�o����窣���Q
�j�cX�fy\�]�\�^��x��g�\�~('�����K�y4Ε1��X^}�t�V��z6���?����7S�ڿ��m]3{��y�|�&��3 Ѷ���T�Z����?\���4!�N׃�f�����������%8�2�.&�ۻQ��r`��OBf��Tg��Ys�O��v�CQ�������w�N��~u��৾b'\�랅2j�	J���p5[��l�4�e��J���<Ig Љ���\u}V|��6�o*�c}����ߛ5>���E4l<ʨ��T��{�����\��������@`��˷�3��ջ,�֌��#��I�|2h��`��h%�4/�r�;:��� PIvY��q���LW�Z��JƋ9�hh���&7���.ȝ=���.nl&P ���־�΅��u!�ٵ�Ic�v3Mɂ��7;�C?�&��t�q�QH%�+�Gɍ
����qy쫺�s��e'��bVn
�9�Wv"�u���v\5Q�(}�L=��q�l�$q�����'��EP��=�B�uS;��u�� (TC�wSە쭄=���`��v�t2w9ݧ!�Z�{B/2Y�&���0d�~�/N�Md�+�,mLk��|�����Hp��XL~�3@ƚؒ[��e�Qt�x�����i[j}�Λ+̪@a>���?	�V��ڵ
i�޳n�ί�`H����0�ŷz�k�{*(���������"h�g���O��<&��=LY~]]y��zB�gsi�%c�oY���~������5&�i�p���7����l���$����R_Ǐ'�z�Ǉ͖z�Nr�l&�6��Ú���ݟc�k�����*4H}]�����n|Δ��W�"��R�^	��\㸱ч]����^�N��'^i>T=�1��`sd�KN�2��,�����E`i�lݲ�PO��\�l@Y�13n��Ta�i�^N�M7$H��:�~Sw��h�>Q�l�o����fpʞ�D;a��q�!ƴ/k������6_&,�R�5��m��H�A�*���J.e�ό�[��'��ѽ�![��=�)�@4L�c^	@�G=v���d��Q�p-�\�\I���\o�'
 �f�譈1��<�ɞ���P�6��Z-�'R�qu�}�p����=̔�V��S��
�,F�	���g��A��)�V��>:{���ϻJL��������'S���-�؀��D�'�ޙI았R��*�R���k"ߛp�TYN�m�ݏ�j͞�|���Z�$���[����X�0|������u�fT��ȩ����TL�u㣯a��(�*龴we|��8+p��܅Ύ��F��N�Z#���_��N�|�vB�
&�]��|�2A���-��R�w�W�"ɵn���z��4�o~�L�u�Teí�4e�4|����uL����X-�/F��PAy�;��qJ����$H�J��x��6�ElR;�#�\�t�E�
*��������!�����=:["�ǩ>Z-�h�i�0KJ�C�y<�V�[���1V]ߣ�7�����>0䳄�)�(�aW�idN�U�쿰�ڛ����GðQ�9�o��(�o�9�sֈ�5au�m�Ӳ�"�w{E��ou8�v���֝����qQ����v�ʉ˭y��_�|�91��ϓ�?wz���`��4ҼL~;�'�ʳ5�oe4�����뛵\�>�H�|�m�ȹ���m0����K����M�pM+!">L�3����:A_X�]w�EFDJb��.��T���A��E���C�����3n�����3=Y�9*6���!tmV���j���	�]�N�QISB�'�Q٤��'������4�����N�|0�DR>�ﰗ�""@�*e=���S�C�#�!Po(��酟6��'�{ۋj�g��(<���A�D8�
{��I�@��I�iaR�E����gq)��������%uU�)���()�&��)�4%Qp��`��J�t��tR&OF8�Q4$����*��=~/��*�t�<�hOȏQ2-��+��k��V����) ��Q��3�%\�V��(S��%�?w����D	1�Q�4+��:G�ewI�<SeO�soz��~*t[F��!a�?L��<�-W\�O*�v��ňLy���;���b�7\�z�gUe�:�z�$4'<*��p��qĲ�v�˼{�s��b���zZ���P�G֧��0б��"|���64��O�A��X���T��dK����`F�&� ��g����_�m�:�h���]��b�jM���fB#�	,)��T��Չ~6�̾�.�e�h���ǀ3���Qn�U�O�(R�1?���ȕs�'fkm�H�����1��6���'-���`|�g�9��ɼ�r]��AB���d��b����|���/?�&��@ )��}x�24��/��o�z@r5�Ҳ'�qjf�P9�6�����>��~�VM`.�z��0��`SE �M.�����ez��y6�^#مċG�#n��^�xՙ`oU`�f�ۅ3��6mF Z���5�w�o"�a���Y��f�iΕ�T��c�A��5�Li!!:��;����(\�?�հ�D`�(��fo�l�L��m�}c�9�����n���mV�ŕ��L�<�<��ok�8*߅�l;%��. %bf\	QE��s�3���8½ǥ��>h}�i-���o��V�eݛ��«Q��#����1m�����d�T���A_�{�@_e�1]+���͘k&�x �xƟ����c��=��a��z�6nhL?��Yx�$y����F��$�5΅���X�3�e�+��N�=��'g�I�.�p���yyj��g����.�s�*R0�rh�}�&�t�-!6�y/�׃J�@	�d`qiv��[�zUaqу<��y"�GW:����y�[%P酔����w�>L��r@zl/�)�bB�͂hO�衲���VT�иu��}�}rjT{�i��pfqQ ��b`[�tF���/���ن�Xpٸ3?R*u��u�׿ V���f�κo����36���>�4!"��gK���o?$�2�|y�F���iv��h m��>唭|y� H\y��U;ܫ��\KY�������iG`UC�A7�5Z]p�}d�H�A$�	���ԍ���/�g\��<Ax�����6���C�Q*z%64i�k�8�Zp��T��z�"��֭-��؄ax�?�# ��03[O����)�C��(��OhV��2���gf���|vig<��jl��ied:	���Qu�_��ɧ�N�t�)�K���q�*�y{z�j*أ��(�7�y�Of��������Vw�Lrq�dka��X��E�l ����L���6���o��ĭh�l����:�65�˸��*ȩl|IK�{*rg/�D7q��=�ݪb�>��䠔�[b��/<\.�궎*�zp��g廇�z6�N�?��*^�emD�'�:�s�]�7s��J|ު�$�hH~ G ?Hk��[�Z���8M��"��&�aۨ�;$�S�
�e���U��օ_�����]�w�ؕˇ7�hf��X]g������N�-�Ц��*	�N��"�E�M��JJ�`����'�r񼨚(�1.��M�#l��{����Dd�/w����Σ>-�<����w���s��q&U���r���<Dh��S�Vr��\�N�J;���K=Ȋ}%�b�T����kv��ת_���C~-ְLq%�6
��j���6����l��R� �y_Q$Z�Q@�4��n@��^pK���X諧�%a�G��s�?;T�+�M�[N���0Ȗů̯���C�tQ����~�	l��x��
P����;��Ւ���k./E`K\��b�?TfQ�+���t*Ɯ�M�|�F0��q��{��*-�9BF��(н9��x���C���.E@߭?W��L�{�F�X�)9d(9�(��<Oo��R���KV�6L*�D�-.�6��ה�%��i���Hh�_Sb�i7�0����E=�#�:�l�Ό�Y�ysͺ�p�d�(��t%���ߓ˛qT_�%����o�gRD">&�e*�E@��Z�?�۱�F����(C�OJ��$��r2n-O��#�_ޚ\* �ad��fPEi�c��7e mm�MI�Y>݁��>���P��i�3P����� D�_����̀=VEN�탲):�o����(�׳��q�}����@8v2�s�C#�GsW�CU���|���ܲ�r����㢜fL�E3EB;K�N�&eX�3��'�'�ׇ!��6��tE^�w\�d2] �|�=r�J,���,\'���IB'�$ڙ���z,}fķ�0F3x T����,<fРl��<��5�ou�+�6������l[��d�1g6�U��n)C	��z� �6շ1���4S��0��n�~U��Ư�l��6�M��D2���~']ڰOAr�}��[�l4^���qw �M�(O`��d�Q��W1G�V�Tb�o��ÚP8�|�鈴d��~�zHR�D9�I�a[� ƤY�z�j��<�9�����Un(�s'α�(�x���P��Y�6����F�4���� 1_���E�'�����0K��$���Vb��Z���Z��R���'oc�*�{���/v�l�1<��g����5�>�u~�WC@��Ё4"<��,J�ӷ��q����V��U`�m�u}�J��!}ۨ��T>�"|�&�"�C��9���#�Mf��`q�Q�'��⏉�?9b�|���UA^K�;z����Ah��i�6M��K������� `�A\���kx��w
ƒ����a߃� #�ߢ�w�%e5����z��KI�$y
B�(]^�3h<R������z�G_=��KS�����޾��'���l������_��دn���X1X&O3u)��2�.Ms���a^��������,Cx�ϸ���R��r'���0�6�{����KɄ�D�uD��9��d-D�e1K�u$��y�K�i��R��xŌ���~�"/�s-O�ʂ�ܲ�S�!K�o��u▘�I����M5�2{ƗTt	��"?#"�R	7;F�H� ��Vg`у���s�	�F����=j6�����7���\�e�"��bF`.&<��5%9Y��R!ʓ� =���8$�2 �2`�|���H�%+	�J�;~'�*l�'��<���]�����@�6��$��������UvZ��3�c�U��<W%���*�r�ɏ�=�v3��33dm�jarN��"��ņY��պYFAµ��Z⩋[�5t�*1룝�q��ڬ�xR�z iqk�Dm��GW���2ԥ+�%rr���담5]���~��f}����l;��6�iޣ�� ^��� ,t-3l�H^��\5����W��R!l���J8��A�:0�pp^n( <T�MD�0�3����"W�8e9��~�5�:�T�$��ߵhn�;b}����{CSxv�j� ���o�M՘�e�_��G�]�$����hI�7Qٺ���tD���|\��x��i�Ư�}&� ��c�w��Yc9�?�$��>�h�4��繭�A2�=�hS��11欮2Qtl;��e�Ya'=�Y�H3� 6�'뤾굑b6+O������l7Y�[������װ��Bqh�&p�V�o�BP�;�#ۆ�+W�E�@؏�&�x��ǈ�dz��[���[�KBz�JA̯�^A�N�!k�e�����e�2�6�*P��/S��2K�Ӿ�[Y*W���T4W���J�(���������-����QE�)�2���a����ZP�C�l�K���8/�*��*3a��H+�eO<��D�$:������⍕�g��\-�s�̹ ��<��k��a����NW���/'�Sbx����;�+^���	�~%�w8GHpO]�l��D�Sfwm�w�P��A��wp;�{�ը�KLܳ��v�@�e��g	k=���H�D���g���B�TB��i�..���΍Iq�
�t]rJ��Z�+I	�^���1��?v�p�"\���A��-w�h�vz4�#ےHQZ��"̲�J0V�)��1[��I�"���!�C�#׆T�o.n�2�=!�����d<�@!�����X=��۫j��������R�S�d�D]�p[4֥O5�F��[s,�>6a�
,�kQ����հ��*�Q�4�����V)"U�v.j$�([��h8I]vu�+���\�t��[����@#��Ϻ���	�+}�L�zv�֦���<5I�i-��/��/Ţ^��|�M����LW5�z�̆��AB��0�P�'Gz�]�~�p������^D�8vܦ9������׺v8np�9��)_ʗ�K�&4��Z��V�!�kJ�=�!L����3B�����P������P�w�(�R��Wλ�9���=T��D+!r�"��Ҩ��r�89����ѩ�E�a�I�&�Ou^�?1?�N\\}W�����̱&��ʔI��.��L�
"M��8�u��,j�~"�\j$�1�7f�	ٟ4�R�6��E�Y�i-
2CP4���-�T�Յw!U���8r�A���\���Gգs"�S���JU�����Q�Ԋ/��6�jMH��k�t������L���}�.ܔ��J�)�v���^r�@:�]vG"U���P �F2q/�bF���ɚ�-� �l��F��\꾠�jr�*���J|S�ZM��ޙ��Y;��;$L�}t�7���$S��K��kg4;i�(�H7d�+	[��7Vlo�<d.�v����Ql!D���L�X�o��.�⸍d"����F��=(� �d�p����@օ��WvR�dh���W����s��̻�Ǡ�c�8�����E,�Φ��B�~R�)	ê���Z�Q]�&��Y��P����Ȟ�^��m,��O���T.g���<9��@�?2��K��5=p�rwC�a��Mk]�������D�iì~eB�%�����������0�����C;K��L�Jx�$󌕯a颔E愢C���i�A�8K���2
&)�̏^Zx
�D'�nQhW�<t�Y?�Z���2���ïH#Ry)�4*�A�)�~���L���u�ޗE:Y�(<2u�ݫ���j�R��%UodU�?���4�o�JUwg�>�`D{�����"���v\�Z�vz^o-�!�	�'�'�1*Z����'S>�q���sw��ЗX�b����9�tY�~�t�K�|"���?�k��ZU\��F��U�L�?֪m@��+�d����$\h�q�3E\�f���O➚;L��ɭ(�UNBy��ح 4�3�r�4p�C^��WL}.07^�$�#W:Q��R�uZ�̕%"UJK�e�^���*;�f�BЌ%�w]�O�����%C(���db�v�"G�R���j�/���_a;���Qz��T���(�+��x@B|�G�#<V
��$��.ZB��k�"��Qw���B�VҧcF.�"V��8�!����hm��r8<Q�v���(����z�m��3��C֮�V�-���w~\�(3Ԑ9�:���ḙ2���0��E����g��T�d�A��*d�3B:r��t~�i�[U��S}��knTd��:�t;��)wA��:'�A�N��/�%D76U{�Z>��`�\��0G��/���}�p�Ѫ�t�M�l����Fn�]n�5Nl��Jm\e�g&����O�^�\�TWE��
L�`=�BY���i@Q�R���+�/J�Ҳ�~O^ y|���������eU*��U?��&�G'L05��6H��r�w�-*J-X����c��'0�v�V�������T~����bԿZ��D���|.�&��t6��O��Gz�5��/R9ڛ���� �����8IW�����f�Y���BM �χbH	9�]�g`���#�>0���h�r����fց�@�ߟ�*�=��c�	ʐC���x������dܜw^0�m"��B�Oa��>����>�'�_I �F��=4���x��ϫwE��=ّZ4�T�ũ����3�������Y�Ù�4OE�/=�c�]"jEG�o�=,��\�W�fH� }��a%+�>M9�.䠏N V�N9R┏Z7\�Jq�:�R#��O��`�������+)�pk�[�����'<a׍Q�����5��\�!�jW5,�<5��:�Xmr\�o��Mu8#M��$�Ţ�T�׸+����Ȗ)e4��6R ���Z�����4��-��}�K�\��[GWX����Za��b+�ו��k���=�g�;>R|��Y���I��lm���N�f ۂM:�D �A�q��sR�2��!�������5ڈ��S���Q?�6=H����`+��T5d�g���oyr���¼/�#q�{DΣ�!A˰�ĝ��N����3	,��vP����ʐ���mB��Q�{K�����F!M�k�|��X�= ��⷗�����(�q���`�Pd~E	�	�qr�Aj��x�F��� I�ڮ���Ą�o��<{�KA@�HIj�B�ZT�6z0�2�[�ߍM�L�h3���o_B.��r�Ob��j��H-,Ssh��/���|�u����5a��,������:ٸ�S�3:̳Z=�,Z��U�4.�Tt��Z��NU���QЍ^VğP���<E��o-}�����6���;i4�Bq�=�{ˏ��:_�"��#U^;^ȃ��j�-O\������	.��4,��%�`�JbP�k2�?�k4�Ŏ��!ʬ���]��}rz�*���؇�'��pi�C��}Qk���v����,��V��Ϗ�y���������#X-�[��QD��u(�E�B��jv�O@����±ޗL�3t�	!mF~@a��I1��Ĝ�>�$]2dɞp�j��]��[<�n�NZR��p����o0-N�n_�4웿D�/3��nZH� M�W���,aP)꿝��Q .�V����"J�t	jBVR�u#�\ʁ��l��s![�ے ��,�����]Sy"�Ԙ�OvI0^�ῐ��ZE�_�T��`j�;W�\Zz�_�N��*e�­d�M(��ve���3O�\�ށĭ�э�U!9��AD?,݅��Q�BsN�V�p��)RL�xĴ�燗��P_g_*�����̸E��������m������y����H�0��@�ML�!K�Y4�P�4�?���d=t����w1��4�^>Q.=�|�,<��q����@�/ ��|;G�
�ͭ��
T!%?Lp�
mj�vp9@�w��?��q6�c8`&������pNĿ o��=��}	��u���^d��q�ۣ}��<4k@�ʷ��>*9�j���h�`Y��`�KJ�Ә�*R�7|������	�X��-�~�
x
:���_8��z@�}C�5�O�Z���U7���]n�8̛k���Q�f�+ �k샯��~�ӑ�jiUQDy�q�h�,���<F6 �A�ϸ�2��/yG�A��ڀYJ�s����c%N��}�:��P��^�pz�k+�0�F��+@T2f��J���Z V��I�����ojӢ^��H�f��>��s�fBX�0�L��m��Y�~�ʮ!�P��|yOK�GQ-Ou���i`3ϲ��7+f�{Ԁ<�)���c�ڂ�j�q���1�@1�C;z�|��iGN��F�P�x��%C������b,�za'49X3?��Y"��%�^�/E7ݶC��7�X�_{���ǯs��na�����R�]ƽ%�����?�G�D'�G�T?�Y6���U2`#{+��p�Ś���+%tߠiO�.��D��Z< "�lZ3�@{�E�!�m�C��)��VLl��6��\K�m�1�_5��կ������ȴJ�Eb	sYv���H�=�&���Yv#[`��X�VwI��Fمd�:�S�+��I�J.�U"[�r�+3�	��m�	<,&������y�K�M뚬�	���>�H�Z���.}^�x�����j�x�����'3����aSK�*RV�G-tn��3�p]?�r���͈�a��R�s�m'�]�e����)x�h� �0q�
�"�V�."�}0�F���>��	�$�����"a5vDAV��-���Z���=PVJ�w5����&��6��&��]H8����b��f�S��i����v���Fg\�Uh�+�_{��	}�h�G�"!p'���뾏���+���Ǿ&.Fߣ���u�'�@/Q��m��7�m���˧<t��7#09���;�Cc�N�X�:0<щ@�DGv����{.l~���|L�d�*=,���l^���tE�Wy<�����3�R��P�HC���"��p�؈6ƈM�>�)g=��h����hI���B�:��Q��#��OiN�^���"���ɮM��(Юt�c6���x����l� ���=�9���]G��M"L�/�f`K ����%��q���<1����u�nT�Xu��z������.��7��r=-�ۚ#� -z�'.H�6k�1+��uN^ﲠ���n���Ц�qحDJ-5�G
�W�7���b�N�/�'O��[JML�[I�96�o�s�⴪�&6Y��mT��7iC�^�C/Q��	�Yh;�
��mWS�����n�;�u�Pr/�Q�+k�I�s��d����p�q���}q�is~��R���Ek �/|�[ԭ�܂2g9�����}�;��_�LI����b�"�Q�hԊA��r> ���c�\{�[��~ߊ�)�`is)�-�&�|�K���Q�{��x�;�����o��;��h�_U;R����"�Lrҗ\|�1�R0�J{1 �4�{6��� y��U�44����F��=�=d;B�K�J}�%$ou�F�rE��)�t�ږ�27Q��������ҧ��B��Bw��L�Iz�!��lj�^�yxl\�{��H��IZpD�%�텺c����$5�!��8��M�IE���s����n�He�,0�`Lg��敉�l84�,|��D7�i��P1�Ch��k6]�}�&�
��M&�<5��G/ G�HKɰG�������7%�`HF�^	N���4O|�ט_$+f�|o:�=���K<�`ֆ5��z�t��Цt3[�m{�+>��C����rj��$�Ȏ9=��l
���&�г�J9����,�LZ.y���K�ޮ%�Y�iX�k��BF,�	11%Уi?���g�
f�-���"�g�!��ql(O�7W�W��j��	�~5)��C,�ʷ}�6��F6wRw􏁍��� �U~譨��b]-'��q&�b���/��e��| k0�`Vu�u
R8w��uh�Hq9{�4�P�j5����5_��C���G�U��n��^(�������@�+vC&��X���`���w>
�nF�et��q��Y��lHb&�{��8���hwsTW�vK:<����T��$3�A�.ǁ���x�x7��F:s!AU��c�I{}��1.�J	�I�E�b�(�`j�$������>��S�s�+�CQ~�]
��7�)j,e����nNn������i┇�ڡ�2�C��d�ӹ�f�1���g�&k�흸	�ꅤ�ety�&��¡bz���"ӽE����3����ٷǼ���83���=��w>�Ş��3�,I���l��������䝘�@w��fk%�����y���D�R������&�w��q��E������v�>?�'�� ���}�n�>��'���lG���2]�|���(��{�:fޡ�6�Xr6�=;��C`Pw۫~� ATkφ8��X'w��ce�2rG&��W��Żð��]\�Sm�B�Ѩ��p���*����`��H�}t�@J۳�E��8����� �i���]k�nj!"��+�	~p���.��F�!�,��<�!�#����셎C��yҺiJ�4����ʡ~�<�sQM�F���lO�U�^�S?��w��0��~�Pf%�81u��N�y֛��rto��h�L�'&,��'�K�e��)3�����r喗�f[�k�U=I
�Շ%�68���w�!
��=`L,�!�O���]Kg㐣�$���������l!UB�N�s'����hv��a"�u����wc�m�mG5��ٺr0wT.���4Jr([��F�<�S����1�5hr��>E9N�'k��N�0vәR�]�:8L�1՝A���(�x�7L��w����
���=��~x���7Li.�D�6N#|<���6�]Z�wI�x��^.�{P�].%*�H=R�%Q��	�b3����C�A����rզ]-Ycd�WT���C�G�WQt�׺`��>�A:Ӻr�3�m�e�Q�����~�	ɺܢ�'�)Р,���u<�:\Rӊ�г�7F�f�"T�.:���J���Q`j�0�p�Q�R����F6�r�0��o�-�ͲX4_���Z.��f��)��ڒN	x�c���p�7�������I�ڟ~5��P����NB�8c���O�H�߾Ƈ�,7����M��ɻr��tK���՚v�%6�#�Tu�����xY�n�n�plx�_��^����wunD�*�@x�$y+���.3ƫ�{"ռoC�/A����]��|��R�x�c�kU����E2kX�`��O��s=�|�{0KS�a'����p|��>�����^�zU�n��:�E�+S_�d�(D�{\�y)��{z{܍f�cD�a�(r�/���@�i��~�X� ^��J/����!DĖ����1}1),>�q�K���5Й��Y����a*/wwI�f���J���t?z_�>�''��R�<�E28Y�aaK[o@�]�p�4c����;!xW}�<�}�aqu�t���c=E����9c�]#�tT���@��������e�kέo����z����K����T��{s���.�B�$l<������0Q�n����U�އ�żյ�,Ŕ�,�伓eM�y��K�3p��%����*�D�.�
k^l�5�`����:�!��ڊ��<{֗��t�
F��W���CQ�]�}���f��p�S�JQ��|M$���8���ī���R���s��6Rm\d������2n��Uu��t�����̓�>j�T��i"f3:�'�k<��y Uߞ��h����-uVZ�����#�Z(�Z`���,�4�� �*����Z�E�|Jئu��U�`��廇�;��6�}���M֨d�
騚OW�Õ�1�RV�`E��_ǣ
�߱Ix�z>.�oV�<UX8N��k�q��K�S���tt�~�|�>��r'?�͘J��y*��
����+��X���I�T��d�*�X.��E��ং���r�$ŇA�6V�5����y��=m9֙�F�H�*O�:m�WP5�:�F�U�� VŶ������<*)9	�SL��&�9\�B��Tg���#;� �^����,���xC�^���˯w�d����ʻ�mYɄ���6�Q��@uS3���Z4��!�{E�Թ���J��_��W%\�2F�ᷓX��9�T�����P��/P�x:�Q�I�y�PP��<���H���+�bノ�J2��zB�AX���֍��HA���Ǒ�ԟh��g|���ܠSn�>r��ED������%��~P���� 8<��F-���b�K��E��=���"/����oa	�{���p,7�@	�l����J];�ܺ�|L��W65<FW � ��@�fn,��U����6�M�ڟ�8��a��ӕ���֚��[�p%�����JP�{_��L�PY=?W��*l��V�MniG6[�W_�T�o��J�T�C�kxT���@��gU� o��[�ua�]@}�o�<�\���e��RN���;���h�g炎cs$s�ƚ�<>�sIo*�קz���e��J�(~VKi�ya�{����4(���s ea�z�f��4����Pa9lo2��ݶ�p��I�X��t����W��!Rŀx`}�-��2�+�D���yG�V�U�d�*V֛���3�����E��c@�ಚ�� ��T�EU
�X����U��$���[�O�>�R6S�t�O��磠	���eXRR��κ�jS�u��l	\E�g�7��ES>%?�?Fk-%]�-�(��T[��Y�����6�֨���J�҈�����ѷ")��w�������' �q
9��R4:�5wF�@ҷӴ���M�U�3v�����#�{q2����2�&���눰+�Ɂ�*�z^��!·�6Z�Q㷨G-
���UK*"�u��g�~����Y'O��<VJ��ɖ���[{Ql�+'�3��ٻ�A����`-
j��)'�l,��n��W���늽&A������oz@�\���5�W��H���k���GU|�BGk�Oh �58���������{������շ�/�!�U-V�4��𳎣�������X�" ��}Z�6�9��������x��E_qcw���8��m�-�����:�V[es�hЛE���̉�p�S_2)�O��1 	Gmw�v���D
�"ȏX,KB�-�&�=X�-��:�)ŧ�o��g�T'p³�uN��\X����⠳q�I���H�p�پj��2T?��7 u�L��=�-x�����0��M�/�=����wic�I���XE���{��:x
�� ��fFi^X��66��l&�Y��vD56_-����,�%��z$��=wm�����8�Ig���L��bk��Uu?�w�M�쮈�b�/n�^k���g�����>��\���S �&��4��<�Cd؛��]5�a6<����@�� ��#����>��Ċi�:_�2.UU���Ŧ*��L)�uR=����F��ؕ�Cɬ�}�jN�f��21�\�C��Y���xxC�)�ͫ�Y���gB�{qr�?����8�	\A:!� ��-�(�J�gP�į[���ً0e�Y�T,�m�� ���B�'W���\)!LtUh<�.pn�Vbـ�/g��ʫ��U3%�X�!��ma�\&P]-7�kf.���r(	g^С�`RlD�?��6�Ao�o6c6\Yi�_�zLW˅6+�I8t���#���w<�#�\e�
�]�0Hr{W������/?a���`pǷw�8y�}�&��{��$����wL�[)�%F��'-*�����U���T��������bR��%>	�������I?��6�be\p +�`�B1�*�dRO�����?���mplx	+�\7C���a,T��:8�i�0G-�-�hd�4��f�2��%3�p�%V�y����㮴���||z�\Q���q�� ����`w�f"��� ���1�4]"��Dx�3���,>�w�\�a>{D����vh����-��a|�����X��%>��ީ��<��TK�ם1N�:��	E��n��_��V>�μ+���`m���{j�������⾡pU���%�b�����������*�<#��Ò�Տ��F9w��Z|l[����s�p�N�A10nA��y>^P���AWL��W�i�o���.�iY�:���j��J�u�
�N��}aA���d)���e:_�WN )�����.�����Ͼ�y��E��PЫ-�)̻�k5�������gp+�A<n򤧩l�5�P�$%��,�8x��?Y~���oXK��67���mS�oX�/��rV������p
 �RO` ������zo��!���B#�NN�ə��;�L2`�ۃ&�I��X�e�O��N�=
F��g(�W�1����>�ѕ�j�c��U����_y����?Xn^66����	iإk
��d�9��;�'�4N���77p�ɩ�-\+*"΄��PGL�����u<D��HLC8��;��ٗJj߯F��,j��mPc^�^�)슧[�͓��y2����w�(�B5�-4����� {^�$�F{vo�'��FM���^6Fe�킱EI_a���=��ekfYQ����q�W~e�X������2�:$�c=J�����"@�o��Z�� �UĒ�T\�9�����OT��~w�bw� �H��HC����n*~9��Ql��JN)?�H}a��ì,�{z5J��/7��)��X�t��Ү�����Z?x�1l������>ȍ��/�}�j �"��Г�Z��Q12�����Wr���,�f��طҳ3��K;�6,����m�{�&q�4ۆ�0��R}c{i���66���\nlE�;�"p_��3޵�����}��m�-|� =��c6���a
\���}��~�'�X��tq@�������֢af�x�<���tva�D��%�����y��߁��P�h�����j�T���Ñ�sS�BYp&$��#џ��U{�c0��e�P)F� �gG��Z����h��J ���JM'�%�	���N.!|�"8G0�m��[e�#��k-V$߁o��WԷ�h5�r�#'��8�>,{��O��N��So��ovܭIO���`���L�iu���J1��yW]f9{!!���
��V��<N�Q�^[Tb��-7	�*ȗ%e#@��2�=�UZ�R�w�w������(_^󁯤���z�p>����ԩ&�#�a��|Gk2;�#vy�@���j ^E�5}2zW��l�\eJUdU��˷��ת0mq����;���x���hN�+��=�L��_�����"-�d����۝D�\�����7Q/�8?����67a����d���[��^N���S�u��.G���P�'I<����n�4 �)&m���G�H���)�E�[�Z�,����ݫ����b/��}F����/sLL��/<��(Ą�����5�ʢ$&�8���N~inm�����e�x�DO����܉{�U���ly��F�썤�{*�3�Sz��gj����B��6X�����,w	)1Rb���>��}���{��@_ɃQ����a��`��bew����[�����j�c��L����~b���4Z���y(� �vW��]���c�˭GvD! �
1���.��y��Ϯ�<~(눪��N�� S�����2h��1ֲ3�mC9�`�W4���)�?9q*8��r}�R�7G)�I�fT��Dx9��dl=C"��f�N��Ӯ�@��2�B��t}�t���9���X%敟�u:Q/DL
;X1�j�(	5?��uM�n�(�ه� O|n���1���H�9�tZ�`>F[��o��K�Fy�Tޭ��nޠ���c\��!�G�1f���6�HI�Z)K(.̪1:]$9���a��H�U�d��,S4�5(e"Z�uwaXV���C�,��;Ӝ 
,����8���I�LT���p{�y�O0tdC����3ߋ�7��,�5v�v��Z(�T�U�͇��\���4_��b	���!��pp�x{��-���J3�Fڃ�6,mYg��Z��b!V�tvХD�c�I�Z�v�a���JO^&���U���^���Iһ�{l͐s� ͬ37ü�'6��$:v�]��������r��^������X&$?���4�:��.륚��R��#�;�r����͂r��J��H���L�m���5{��9�I��`��bX�U��������yp��\�
�*R��jQsg���؄�F�r��o�i�:�5E �!��,��p�
gq��dT�;�?�q���ŀwv( T�|R��Ҙ"�m^h0oU��d "� �j��{>z7<#6( 6
%�p�Ư� ��OI�+�����zl�ʋ_�U���i���>էH)�.EZ�kv
��g�)���vK�h!�B��u5Togbe�LQ[8�����x<貽�{=�y5��%%2�5K 1�	�ɻ͖����cl6��[F��ߪ ��sIU�*�0|v"q�G(9�ߚ���+�Z����=����yk4��$��
m�WnY�EK��=��M�n�Dg8^��W�y������3~;��ӪCRи4��0�Lo�55�U/ �)l��d!ma��w�/��H�;`�8�*'������(9!a�y��j���u}�1�֣�Wm-E�p�`�%���
	�7E�	u��)mU��� ދ#ABRK�e܏'�ġ�Z�ԿP�/kw37(��J��_o�5����~r�du�a2?�����V��Ƣ�vu�`�F,�s��j��g	⯈"�[M�a����(�y�Vz��X{f����m�
�f?�X%��iL���EWQ}3[1Y3h�������s�N�X�\ 9m/.kY1��3c�OK(Q���@���L�=�ޝ��mՃ!*I�H��ծ������z`�;O�y���´Յ�7�����@CtK����m�*�4c��#�q �tO�F|n�jW r��b��hWt�ad�w(N�(:�4^ߏA��o4v�T�%�� nS��׊:�1��&x��HJ��uX����7_�L��-\�NH�6�\.�����v�߀�<0�(���]�^��;w��d
r�F���+^M��k4��h�kaH������9�
��R3�-uR�dq0?L��c�2U�E3��N,� 
_麅�CUx�������y�#TIɌ���Rɽ�����8-�}���2�`�ߨP��m1����(�k}n�)��שھ���b����>�r��z�4�s�",gz	�P�g_B�c$wh�9�5������>D���X�@Y}�$�����uX�J�Dw��$].
/��=h᫑qu�<�l�,����Ȳ��.��r)8.6:��(�؉0��dh$� ��@C��B�[�7��2�7k؋,%:��퓞��Q��1v1�ę_Ң��%K�{pS��{���!~��a#�#W�ϑOKC<�q	�F
$�#T̜t�6��S܃��V�Ma�1�Z�褌�͚�}�SR��,O�2i䪋�"��'ʉ�ߔZ~~����޸�/���ǿ��~�۷�i�R	ľR6Y���#��V�|���)�Ǖ3�E��4���if{	쬊�����+�W��l�
�a��*�c{������������%��Wb�ߠ}UΖ�3K)������R{��37�n����/y�����Ǒ�m�j�"�p�u�B?3��ލ���η��n��23�u��v �+KYY&k��ꩳ؅k],cK4�o���ï[9��k���z��c���*���`f(D����
�p,.x�w�Ȳ����D���*L�5�0�u�W��i?Ka%�sB>ǡ�����72\^�gh5����}�J���~�R:�Ϸ�Y�t��K\Ecդ�MZW���ߝ�������p�'��+��V��$�Ydۮ���F�q��\E�L����^���OC���u��Ĭ��#@Q'�T�N��ṘaS|0��+N��>���ѓ�|3n�cSU�7��"D��~���<F�iA�wB6���(��m_�)2	˧W�u=	�#	2IÇ#L��E �@�s�=��׼��+����V,�n�����t��p���OR�:�k"93r�Eh�}?�wIc��^3�'�#(�}j�}�t����ҭsO�2� *��c��2%�2<�~5���a7�+g=�;&�ic��O�Wce�3ż̝���d6B8?=l0Z_N��?�*�?��u�L-6BB.]t�E���I��B�'l<2w�)�-:�U��x����$G��t+�*��-�~����Q���:�7v������PD��*jÿ���K�|M�%G���o���>�����q�j��[r�颎�q��R����E(��f#"�w�fiK~Z���1۲	�n��'ʙȂ!pԳф�1�䢊�Z��nrh$P���_"S��kE��P�/͋nѹ5��Mre��G�M粄��A<N����?��э�ӿ��Y�Y��(�=�m�i؋_��i�).sl��n�����Ƈ�Xr���NR=|��g�̴^y�tH�{Z��
*C��.�]/*��|����^4t������f�tP�Eh��wT³\}�nD�t��z�h�]R7�w�"��N~��!T�Du1mM��XN�� �/�ȩ���cr��2�5�	���D�I3�8A0�֡u�]/�S43�3�
/�410����	C��C����ض
���UF���N9�Y�������_*�i>���cs�볘\H?#���wF���:�RlӋ_�+�o���,�ງ�DE�668]Ȃf
M>!�*�6A}�����N���;�|F2D�9�a[��k`_�#p���H:+}}��,��C��si��*�w��2X3;��ϴ�ذ�@���w����	�����4���ݒl<*\n�i$���ϟ�K�D*��͍�ڕ(HŰ�2�#p>g }�2:r�ã?��=�i�5 �c)n�&ч*"���cN,�������e�qd�x��`.��?2��k�m��
Im�27�)̷��+I/�o�|���e�;X��M:m�c�8+m�̃��� !:�{7bE����QS���K�u�Y�)�ؽ
�$ �>}�w��p7V�����^��j���|�ӱ���YA�H2H��SmP>��Mu#�&�桠u�GW��E1�G�b�%� du%�so7�_,���%��4� @��:lF^��n�D>]L��7q�]�c#$z���h�E17
n�u8��Zo���B���l
7���c�w���T@-���5W���\��d��ۑ`R�Mb��>�mk��3T�F��0	�Ul�mÉO��bvi�+ɬiR@��b��:Md�����ݍ��R$s+_�Q]�T��P�w��8����C��O�A�d�LՈ%4O���n}�h8�.I̺m=�f�vtm��ҹ���dΨ�k� ���J����S&�[b�H��M��Lr�;�y�2]���YH��F�c����%̜�\
��
d��l1����eъyt��}7l�Ǔ2w>Q���I��;�ׅ��:^vk�,|�
P��Ah�v����9t�j�B��'Tɮ���W7��Y�9�R�����y3�3y��V污^&�ت(��>�%�����z>�V7�Sz��-�[U;jՔ��zy��C3}d�N��PL+��I�	�>|EW�9�;
�@��;d'Vd	�@��i�5��1�]K�PYFT5��^��!������mH�i�%��A�[M�M�=�p
��Dh�"5{'�E"8߱|�Q�]��z\�6��6����Ľ�̖�]j4#���~'��&��?L�|h��QP�����&�������ҙ��h��)&�{��$�g[qk6N��2J�9�s%9B�3z�h�2�Z�J��>�T
���F!��49��y�Y�t*�p���=�`,*� W�<�8�4�n����g��ښ@�ҪsՄ����Nӹ�%�Y��ӑ ���m��ΗW��������=�S��8��k�?�Qʰz�L����V�����ų�B�����qhPr|�fL�yN)f��-w�Ap[�%�:*�yk��fTh�H	ɍ� cT�\����
�c��8��p�ZzA��}OO��p.*e�d�HstZ��=���}�)ݟ�Co �D��i_�R'�s_G��hc��v�J��XV�=��Z��(�����K�Zw��nz�92��ii��H����U�,�b>⥄w�����J�ڍ6i�6x�l���!@; �+UZ��Uap���Cn�����F�~DJ�ǟ�8F�rB�xxtt.�x�u��FH��<5��3)�SZ�ݬi��������y�,��d����B�8��<�O��L�xǞM�;�r�$du�թγ�O?
�]��8��HD��Jf��"7Сw�������R�\�a���r�i�e����9�����������0#=�я��?-��sI�b�YC{�O�̈^���+���_�@]��p��b�u����-��B�p.�SrgP���9/�mks��I�.���K�����s���k19��;w�I�0��}��Ӷ1_���It�/>�Ri,�O5����7�WN �S��@�A3}w�_Y�W���K�Ϩ�I�o��f�ѯ�%k���Б��ғ����:��Ν�`RFأ��Q�>L�{a��m�� �k�?v������
�h/��*Ñ�g�[�X����f����0�b� \|dqp�����3@k��d���"�m\ɔ;C݁,��h������ԏ�	4��ζbN����xw$yY�W(n��%��^Ȏ��_؂�;S.Ӱ��ԴK8��̲]�7���_'^���}�A��䣾���:��Ug77ڏ_����U.�3dTX.��]��W#]�>�]j�ZM���y)�]	�W�8
��r��Ԫ�={4�A���G�dSC~�!w��ѪE�����.�}ĽdY][�����+%�sn�v���!<6$��d�ϫ@� ��9!� ��Vd[*<��!lI.��Rdu;����'�^'9+�|w#=%i�� �)��3�dX�L�(�Ni��ʮ�=t���(�qS��%������)I���j穠r_��x��M٘�uA�ӌ,[��½�_�g�ћWz��	3k	hE�W��R*�.��^W2���jsu,��\��t��#,����C�F�d.�Zo2!��\�/����L�0�
 ^�C�1�1�0��>`s�"��z��GP��_<�#l���L�:o�s��c��r�&���pz0ܯ��fz�Y���`�c��e�w�{�3sj���vf�e�GNy��Tb_�G�Je(B&?�s!���*>����g(�#B�E�P:��}-qQ��O�]C�B���;]�7R%'���xٍ��I�$ܴ�1�����Ao|���{~�p�m~���(յ���"�ʚ�]���Y;��*	�vb�˞����F���7�Ov'ɊZ/�Mv�i̔~�w�g�L5+���Ƚ#���@�}��=e��������U���[��@rq�O*?V�l4D�����Ū��_^ *	?�C��/q��]]�>9��'X��T2N���)5i\F��X=��L�I���&�r���}��(m&����IY䒕jr��d�,�T�~�����2�c��x�Fg���[f���'aE�� ���
փw�A9�$y��3[�?��^�N�5Cw4�����oOf��t��G�Ԗ%}�׵�����l^	����i��Q�~�΋=�UX͔'W���1�����n6�#�*KnIf-TZ3
�Zo/M�OB�tW�G�*���k�p+�����>�/WכH�NF����#�5�����R7��9��yW�����%C���gũw�ՒT0� ��6K���$�K��PJz*�{�X�����!L�4� ������,��"�Kc9�4E׵q���}o��bxň�iV|Y�l>���}�Nz�U���ID�S%�-CH�:�A��f�SE��ϩCjy?N���9E8J2��a�5su�L^���lɼC�{�%�t!��N�J�.:$2nlN8����R�_aD�������>p����߽�@@w�r%�f�7K�V7�Y�F�t�$�	�ٶ�w��1P�����*X|	�����&ʭn��$���椢W�#��a�sR�jN�>S�w`��W�A�S-H��V������gYI�=��D�.�&��e��<t5DyZ��.X
P�d,��?��f��1�3[Q� i�6�d��hD �e�4�6�}�!� �x��9�F��$���?ܴ;rCA�*�E�k筴L�E��'����!�^O��}�=��� ��%�L��3бZ��-�?0�I�!��)�(�/dQ������cE�
�\s'�Yf�e�wU��4WF<�8;�5����S���H��N16���D�s�d�w����b��Ȫ�7s<�<Ш���WxD��J)�Ҫ2�E���+�XP��{�@�,zш��^������2�R���0{��{�V?gͥ���g#%�$��ku$��j�C�s@{��/�-{�1
ĥ}35�w!CI�&R���x���9��Z��)�t�.��$�b?���@dJ�� )�,�&eu��z!�2��;�>/����0aG߄� �UJ(����n7\#	�Ԥ���%�t����9��
�[�������pԧ��3�w2��r��N[����Ȣd��s�"I��ٻt��93jH�'Yj�tduo�)>�̚����Tht3��$(6���jHd);hm\�YH"�@�{��],��(�b8u�^l�ƕ]^y;`�o��wi� �Xy�
e<NC����ǔY���P4ZMSR�P�W��4ؚ6o�:�������H�Y�W�!����EX1���yl�:��
!���:�
�(%+��nK���P���*t
JΚ��=�|Sii�Y��[r"9U������i��yB��]��c�3����׸�w8�˳�$m��� iXQ�!��h�N��3Q�Z�HlL�e������"��i��f�+��|��� ��W��"KW�ז|�_�Xe�&�q��ƥ0���b]+*� �n5���%AG��1ԲC���[8DZꄆ.P�9b�:S:2��cà�:�uKk����"4dr�|��1.�ԗ��֌@�L0�NN��PPm�.2��<@lO��=R:�$l�OO/#�+�®��u@�Q�-Z怉�Koר4�z���>�䤽�cF��
�0D7�Ͷ7�7�	˒|�Q��6lܐ�J$����椰:�U9�3-X3�V�����s�
K��?��i��0�o�����2��Ď��n�|{�n%�A�l:�N/�FRJ��`;�4y+a�L��q_����+���+y�AJ�y>��C��Z����Ģbg�#Ր~����owΒ�x�qT�{��U�^��%�:t�	ӈ?�������+,���Ι�l��Z��%<*��U^ h�=w�����wd��6�R����Ck��r �D��5���Sk5�%��áـ�	Ɣ���[��&�Y��l��U� |��9�����2g>�-�]_m`6���I�G�8������*ٟ��a�f��%l�����[1,\l��IʘD��Q0��$r;�?�E�Y�T��6�NdL��sq�q4yһu�~)��.lGӍy��XNM�;���: ���48۱F��X�dE�����P`z\Pg��~*Q���n�ڍ��⺣E���0��$hƾč��dNz8�h�o��(b�le��pV�r��
N�):F�ٹ̈́J{}Oc.72�jR��q���ߔ����$���Y���}j�a0�!Ӎ]�@<:�c�:zA�]px�1�����4*��`o�Z�f��'Q�m���^���\0�B�o��q�ӟ�u����ȨˡT0�ޠ��5G��N��MG W�p���������+#Q��v��h�����ه6���a+1���a�ʬj��>k�֗�x�̵]�qQ�ԃ��A�o���qPH����~��todg��_K"��^��h.��#�s�C�׍X���I�ݟ;�tvL�m	�'�<��3�g��ƮY�BS��n�	��hoc��y��m�SʥF�NO�;o���,-e0�	�:���u%�n�/W
�z��G�ֆ41���o|�����l2�����J�W�{1w9E�v�M�Qp8��t��l��3O}�������x]s(҅�n�����?W������ڿmA�<�
�x���k'����ǝ3�f��,�cy#���(�s��y�*1�L����$�α)��z£�j/t��(eb��$���S�\,.�a�gE ~1�b��>�BI�f2%����Y����&� &:1����O��
�>��A�$���I����N��]�R(��˻��I]�Dq~c��G"�� ʈ�'�5��=�1�+�5�q�v�t@9fg�N>��(���K�(�- �i�L�HT�w_��:����J�a`dnOT�^�&�|FBt��{em@��ûA.g������Q�q&y/��J$�+Z{��rV~��O'�l�\Xh?�����v�bW
j���i�+[}�>!,�6f���~˕%4ʢ�����7s3���#�b���b�ag�|�LW��/K����褛�=)�1-�ǉ�[<�0`�a[��Ѷ�Je���Vb�%�n���`h*�g�z�~uXo�ځ�]������rը��Tt-��1���Pv�t����V��?��J��[څ�ҮFN���ݹ*���H#�����>P,Q?��^�t	w��9�MLW.� �ݧ�aK	��L�9������O�� ��}�U����F��}�P�h7r'��_�Eǥ��8��@9`:1$�2�c�Jf!HLd)֏�����q�.��>S�U��=K��gTe����"��<�������?O�rwjr|����g�7�?d�6�e��%V�g/��8K2��8��!z�
1G������v�����NG�i�B��K/kr@����,��t�I��<�,t�K��[���G��5��׺��zPX�M|�t�
,�wrxm�[Q�=��d����4�Վ���
���'/����C��_/G!V�N��Q����c�h�mt�u7dӇͩ @�+B�m�sBIYND��V#u���{��X�Sn���)��LD���8�e�0�חr�(�������9p�1�U@ڡ�qM��Q�e�����OQ���)�ޫ����?����@w����|]��U�Q`+�We��jR�P����Sk��]������s�GHVѦ�wt#���F+7�"�⪯�t�6W��
�K�{)��{{f�����i:U�U���{*�]#M�c�|"��{�i���!�n,Iڏp�`&ؤժfb4��&T�DW���tv"�}��^���lc�I��J�2�9�&���}ֱ�+�{����;o�M�rV��@�������[@�ڻ�&����<��"?ڨU��������r���7jw���!g����}��+�N���4�����/���~�JЧYc��,����AL���B.0��O4f���m/-�nr!!��c�e�֗�w�D�y츚j@�c��PWЃ�y#��"'�}��|����~(���T|d�ߛ��&�'���JG!U�x(v������� U�
���x=t$����A�Y��^I�OlU�J�z��U�(0�̒>|�BU��䴩S���ғ����'}��
������\���}7���T���.��$�`�W�G�\w�Z2��ݫ��2����(p&�b�ؐˑW�o�-��Y\{��쬼}�z���W�NDgh,�9���z����f��r��eI!��N=����D���/��G��l�:b+!GRα�|3��ɼ_��?K���X���{�QP�G�Y�:)[;G\����gEӇ�G���ttI��*�f�D5�Oqx��G{D�㊳�ͷ&X}1�>�mc��M%�8��𢔅%2#xN�p~��F�!u���wE���m%�3'8��T���`�Sk5���W���Bz>�{Is����R?��[UA�{��� �3��|Nv7z���>�3y��y�Q�/,���������X��5\b��*@1�L'}�8�ؕ�2�iܢP�,�^/��pw��U伒-s���� �Z�-h�3���u��~"͟۴>�{��2�T��+�����R�T楻`�-Ϻ�U�g2�o�T��]ڊ�
iɞ�Y?�bp�8�~#/�)���y�����Ӧ|�Q���.��'.1�9Q��n������I� �6!�O�f�ೇ9��׏���E�Ȣ	&|�����Ņۈ������rC�-#��F�g�'��2 犜���-/s��Ɩ2��	�y�e>�쁵q��S�U��zaF�J��~��"���<d�+S5���;���R&���������:�@"����K�;��'�����5 �����|V��ZBB���V��.m�з��;&��&��$}!��k3f�}����Q�6�=z��M�{��m#�(Ay�2�'�����LlO���U����8|?�^�k�@��u-��� �D�6z}��'�L��Pٓ�B`y ��o/�`��_G�z���?�7��I���aY�Vn�^��	Y�@i� �X5-�����4�����h�����G6Wsi� �kt>�n�J�G�*��Q����=��k�5Á?o��'8�?n���B5c9�.��!F'Մ�YGI��m��{�dI�}a�=�����б'�g�ob�'g �}u`�?���	��������oy�G��өy��j�`����gy�A�o��؇M�I��#.��x�^�v=�`nfp]^�~�q�V�r�j-��I+|!���LDeE��O�(�-X�{!1����͙�?����]������j>N�>rPf��I�+���J�YR���\�h�4�$J�Ŕ V^$&nc8��1��n���m�n�!���Gu�h����i_z�#7�5��C�i�ɫ�Nɕ�9�.o�b����Z�`��1����N�m�ݛ	�i#ժQ�ס���|o SA��$��s3n�����8ݤ�!�f��x�;�+�<�����I����pZz�C;m�s,$b�U��x�T�t��!�:KȈ�]Z���; YE<�_��%]��j$ܶl7�$`��N|�� �V�jp�e[�!Ԡ��݅�DO�+�/&��"�z�)^	�*F�9�~~,i��=CB�_�+I�'�TN�7�
�m?����VN`/���f����?�f�.��p��t�)�"d \�0"4�Ɔ���PW4G0Xd�3�q1�M7�����AI��F�虜��4�L�U�˝���P�gk���E�O�y�ұ���\c)�x\���&���7m%	"��e�3��Õ�_]�ϳ�]�VT=
��w�)HbZPwjܖZA�B����컉2�]G0O.f������)>(�Ejj4=Q��6�)�w2S)��h�㙤��#V���4m�ꏨ����M|r��P�2����W	Eߌ/��ig��8#�>g�W��B��
d�ф��&-B�������Z�O��q�kWE����9U�E����Zvu�QC�R?B�עz�\������F)Y��,�H���~�8@�h�2�o�qW������R��5ƦV� �}T^$�4(੹��\-S��VsF�	�W���k��s�#��L5(��_U2ըZ.�,�m��7�*��1��R:l� �s4~����C@�5V�.0��g�-:�M��=�����4�c_��!3�8%�̞� �u��7M�e&E��};B�\
/�(Z-I<�1P ~�W���ŉ*��j		��g�,wۂQO����ފ�0����������C!��
�ã~������|�t�ۦݓ4�?�2نH��lNN�gl>��<y�:��0�A�@�*��z�������g��!������0�z1ʺ~��1��}?�/��R�{_�34-�x	��CG;���Q��pg�m������A*�˺z�DOAF���~>g�����CC�9�s����q���H��JP�2���o�ry�>Iĸ�N`��n+[ʨ��&m�؞�?p{�}�d'��x�)���v6e�aU�*�(Sx(���[~{�O?�5Ǚ�bl�#n������r^~��%��|;X����E/(����<�읖�m/�[J���h���8DNÙ���1j�R]c*���|�Wi�@�7�����[��#����oN��4����?	;Lo2L���:�%���m
�/�����³3��3 ��QQm6�B��Cz|ݗ�Vck�[U#�o��g�1j�x�f�x�&r��u6��Jt�	���s̏��x֟�W^� 2Z�.�:�N�$A?y-�t�����z��-F��ޏSR�S��6���/q��O�4�����n�i%9�I!�Dz6{�xyG?�����@v9����Z� p�bL�*n��@.��?煽��;�Lz��_����kv�U9�	�~&�y�����Us|M	QN1\�e����3H����U����I�*��	  �blX���*�H��T\|�4�.K�6���<���a�ٴ�W�0�9B���ȫ��J0��+k�n>_Wf�Fs�|�6�h������P�r|���2�( #�+�|d�B�J�1?�ɽA����L����4f��o�'i>M �D��T3nݬ�ݦ�2��-�� 2��|lOj�/��]��7�G����y����s�R'7�$-���Q)1UB���L]�.n�
�]?�.'+'ʗ���� N1A���`����{����'��W2)9(^�8�6��Z��{o�U_M��IN�B������.11���W��AO��o��?��ľxGg����?f�H��o�>��-����F}�l��P�aؔj7ǚ��|R��B��ר���E,��'��YP���z����x +�qx&��BZ6>؅c%~U~���b�M�[���ds0q޾��1B[�+v,����]7�z��ִ�IsSY��òGްʲ�tBMݗ
z���s��iY��H�~���=Kw\q���b��ZX��;�������6���ӽ��\ϯ�@C=-yΖN!��0�D���Θ��D����<&vːcS ���iO�cT��N��ڥR�Ae]��BB{ٿ;��d����]xrf��~�#O�^A��kT��t�C=��w���y��ɑK��M��!R1W�[}�+6���:;�8s㓮���\d	���8Jc`���S��J�������|�l~��{?��F�4u됧=��$�
�?�&��V5�?��E4_��6<f�M�8��E�K�&`[2Hڀ�Gxy��6�)8�:acr���!f0ig��)t�t��m4��fZ0sF]���i�������4��������[��ݶ]���+i�QJ�(:ڤl��%�[Cx9�0���TJf�e�<z�T�����xF�Q���!Gj�^�1��9Ð-D��2�'U*�"!�� q4f�ժ��Q.P��C�YqcƑ���j����Bk�G��cca^�
���u��S�i�n�l�i�B��l�N�%]�ԗp\�Qm�jC��`����I����� �}i;�0��R�m`9<4��N&�p�-&d��3�W���iQ�_�l��,Quw��q:��Y����c��4ER�,�j��u��r�2o�}U���� ��Y�}ru�����(Y��q�u��$��"o1,�s(�R��ւ�]ޏ�k�B^t�Ǝ�\NxN�����������d��A'IY��JT�8�E;x���̘Y4���������y2:�SeH���yM?{�.��M�G�X^�*f����F�ވ�����EՀO%eC9`�&���4��6h��g�K�p����G����I	T��-�Xvn�m}�t}q6;��3h	���E)��%_H%XU/���I�I�4�~�aCs#Tj�&v(<0O�$�c�����n��heB��;$�	9`�Hಇ3U�+�G��I���'f�WҞ�K2��kXT�Y<����;w�&DKIh��A;p����;��2iG��Z���;E���v���H��3��I���d|A�<���D3�0C3M�zWEHd�jU��$T]7%87����.]�R�[m�����ב�e�7a#�㬻��ܫ�̍j���O*���n�i��$EIf�A͝D���7��@�s��}6ඎ��s5
��G���0%�\1a�pNq�=Z���_�t]�rg�H<�ꛈ�"�9tGRBdSE�opFd�ub�m#7��Wq�N,H�;�No�4�$��<_��H�"��}�*����S�%�;6�
�'fJ�:���sp93z4Y�mkB�,W���1��^�� �R��\��2N�U@�������E���Pc�I�J 0Fc� W�Ħc7O�]���ϫ{>��5��J&GV��ğ�nmx;�}o���e6h�Z/'�8�X�}g�#�8���q�""j/�_J��1������h��	��Pr��]G"mn�Ik�ܞTv�G�$�1�]P��ËĘ��)|���{T�����b'e�Lt(���k�\����ī2��mo�q�pQǕo/�"�Yg������P�	�IX���Fow!v4�ۤn�a�H>M����"��r$����*#�w�Zw����P�~{ec-��٦hb�[<%d�P@��i7�2<ʫ�/;�L����Q(o�uH*&��	'y����~1�(�W�+ R �Ȕ�nW-x�qi}w���;Ҷ��Q W����.���i��j��pV�95�(a�8h?Ő`�T_
�ޠ���O6�j9�Lg�)<ќ '�J�dM���nc2�e��X[�$�$ΦI=/[G��7n���,�P�;(Q� �yd�#�3�B�:�Գ�d<�c���5tR�z�`B���e��S���?&�[�6�j2Me�Ϗ
"\
�Ih�{������dZ@L0�+��\�F��5}w�:�1��B�t����	T�Q@�'>Ch2�e/D6�q��Y��;O�2_B��.}�O�%��dd�����N�b�����B��|�vGS,��#���vlh��w����L��g��,�<�N�r�yMe܄V�A�Als/��9�{rv.��}=U�����J�~�y�#����?��.�g�_�b�0�Hbͨ	皭��t:/��åK� }&��b�}�����H�B�=W��#&��6G�Yw�Z����Zm��j���8�X�_�h��h�����k�����v��z��I�#����}�$JV7`���㙍%?yhJ��A�q� �&M��,�.���N@�*ު���Z��h�<W��E��3���9%���у�+tBft �ݔ&bP:��b��q��`9�0�{Zt�P*0]�g�����놯1r�Z!��;��?����"���d�߇vl|�/x���dB��\��H��M���0�8D���ug�, �e��٭���Cl��lG,rDv_��5S��TS>�Nx�S������%��.���W���9yq�އ�W�RT�A,�{ !�X<������E9�$X+����>��$�2���!����(�vNw	S�&�N�v�/%�-#P���Ixk��`q��0h���[=��~_�c�(Y��z�B�gь'�G�W����?� �*h�Ț_ ��jW��{���F�@�҈m���*(~����fM����Xz�9Ac��C	�E�@WΤm@���\Qk��QL�/0���t�c�Jc	���2/O�3c��2|�MTv���FB�~Ո�E:w���C�U�N+��<N�*�D{ٙ�E� ?��<��nd��&���:�%݋wbrg6B^�����ϔ[yc`�$�q�e.��fsD??	/��7�)���S��W�窏H�����$ڀ��9H+`vA���$ˌxcIp�U[w: ��7�ܺH��?���X��qpe^��A]�p���$q�<�Z|����a�]�u6 dh�kü�"^As8�L������BP���H�^彋���/~䑟���$:a�v70iHm��h�n��VN�	#d�E�sy�̈́�?�Y�uS��)&�H��䪉L��.	�U[�il�݇���-ѐ�s��*4N�]+�~�P��5uu~�|!a��a����T��Ia��UjB�_S�clc�J��~d���)�Q�?8��6i{<��e@�
̗1+��[,����ve��,�u�t1�i�qfu�}�O�~&���Ni�}ր�3K7�"����D4�$"mZٖ/��Yz�i�R��*�<���L_�����)����7	��Xnw�> <.m��_�<�!�.CDPÕ8�ݴ �)�:��£cFn�q�6yU[�`�{�=Օ�J��2�Y�m��<��D��^~4�����%���)�����������K5�TV&#��}_�do�gQ"��%ώ%��yv���d��b��I�_uة�`C�z�C�BT˾�� �~�����ad�d�곾����&j\dN�ꇮ�d�	^T(g�_G�[�{/!��R��c�|cV/�t�	;O���$��͙�D����y9L����,�d9��@�N���X�P��Js�W
��QMHߐI�B�H���7KXK�?0d
M�����ymږ�>Wñ9��J��cba��2fl��NB���\jI=x(
s#��k)7��@Q������?��զ�K̿/�;���5��M�0h@��5��K��b���7�� �{f�\d�7L1���H��z���Ȋ��Ʒ����;�E�댵�S��fϋd��7H���' ?�CG˸h!$�q ������]~��DN�w%�/�'O
�����T���+�7�*Ls��b�S֩}#�<?�'�y�"�'���T�Nѓ�F�������P+c�����R)N�9�fQ�ۏ)e0����Tp��tJ"�Q��Ap�ҙ=��6!m����4MrƜ��O�TKCn���@:�?�3�i;����&	P8�~���qxc��Q����·Y�G�u��wr�� (�(�{co& ��!O�S���3%��mިqGàh`!qlO6vd��	wS��d���pc}�m�Yޑ!,��<�d����t����<�G(ay���#��g�oQ.n�y*��YRkx�2�fBkP����^�~��S	,�"�A;�Jr<��᛭���;�_�̃��W�y0�Bӑ�j�y}<�"�+v+b�h�w�xn:Yq����v�6��`��)�97tӷ2��Nm�
r�'\�8O��1�}iîG��+	�c����A���9�'����9�-I��� qe��䒲 �����Ys����,+���[�F6Ϙr�0Li�L~��j*�����Z��Cr�:�=4�`Qx�1M8���e��� L���S�����i$����53�h�n�2�sOLLI`�34a�R�_>��L^�y	)@����Ւ�8��e��u�3 r+PF`��&��<7�0�%��cY��{5�k�b�b1EŘ�5���}o6&��j��'0�?���i�˹���U���5P+&�К���]��<���F߻�*I�*�xt��g�k;��u��H�
���H��ंeu^�������aѷ��~x=s"�'�)L���Ta&,�:�qM�V>Ճ?�*�$	���# @�	&��Z���jQ��Uov���������iG�Jm4��4qЃ�(�~&�o��1 ���|btILŪ(��)
��9����o���0
��AD;�_�E���<��]��w�k��g��V��h��hgҧBgJ��E�W�;��ژ*3�1%���J��{�̬0����KѰ=�!-t^XZ��H��q��{I��Ssۼ�ip&^���:o���G�a4j4�ڴh������q�9-r(���D'��'s�q�_�lP������w:l���olu&�>RWr�z�9� �ZE|�����r�K�Dh�����c>Kg�Ŗ����jh��U���~+b�<��]Q�5�k+Ý�T�jU��[h�|5��א���7TTe�#�v	FF/���%&f��^[����޹�y��ț��|�J�V�+
�J=U��[�T<�#œAO�!��Q˒�Z��u^��}&�"��Zhp��=��}-�&�G/t�w%�G��[�����ȍ���<��\Q�6�ϟ{4��_����^��8�I0����d͑%;��"��3�pB�k�����F��\�f����fgQGV��H�%*<�^[���(�`��h���N��M�ƍ��!˻���|�����@��wu|�he[����˝��n��5��^�Q���jh&su)|�ưE��X�L�7W�h^�r������*bD�]E��JѬA�sZŷ%!������ۉ�Z�8z��秇3��p��Z�)���$���ة/|nE��xN�5��sZ��퍡%#��L��H�/'	�m2�q����+CE����"��wߌ]<�kh>���g���gKTd}�#��H�6F_nB����������Zܾ�+ͩ�q��ݣ̫��,��o
��(�D����%�v��k�?7�����u40[ ��'��r�ڈ3��Qkf����~��4���ͩ�?�G�?��A���HL겶�b�v���@�m�H�{nA�������V�\����;,��m5�e.�w����r,��IL���ڤ����c�N�X�ςg���r�wb����� �SCy�蠎��ҋ}��z�A��c��=�mq9.5��r�	�&�#���LP��AU�o���[S�L�;>t�W�i��}�𓕅��ɡ����F��A .����x����M�G�1Mt�PV4c��	�F0G��Il
|�ٌ�΢���$���.e�Nv�s9�$3�f��7	E�Pk� ���L����YG�w���ros�tRk�"<Lr`+�z�Y�øZ�t�؛Y�	��,����QE��K�I�q��{=��մ��۲8(1�B"�#��9m�~����e��� P�~��^-���0�Iã*r)��l���Y���(���B�o��ʆ��]9�����ǘ���%��?[��p�v����=oz���m:��5�j3�pc�J9�V��V%E�U6$���̒2�XJ`	�_U��T��������Z�:�7qpng��m�f���_�,����.@~N��9ys�M1s��6��e��յ�\��`���^i�A�xV�#����ƒ;�2�Q��� �v�9��{0O�\hު��[�i�y�]wP=ȶ�		���������-�re�s�ut<.>��돟�ӧn��7~�,G��oŹ��U�X������\5v��~�x����8<��e.H��xy�A{�O�+ȩj���Y��bN���}�˃�~���~p9
�F8w]/��Q�Yzc��g�����y@��Iy+X�Ҡ;�7�/B�\P�3��h�d�xP#s5�� Ԉ��*��~~V^ۏ+���������2��y?�����)�RZ�iR���Lg-{��K��s\��4Q6lUթZ~<g�>�8�!�/��!.������J��a�
�¯@6�Em��u����D:h�́������;{+��6<?�y�j��uf�8�b\�P>u���s�%�*��	�c����Mi�Le90�;��kf�$+�������5�K*�4�᯹���� ��@�E8K��B���1�a�鹞Q���s���COR�Zk�����y��xf�z�ލ�l��j}�M���o�~k'�w����Ӎ�@E���=�Б�����4��F��e���cnRS���D�p���Y��
�I0�)��בtM(���,*xm.LxR�Tr���9o����].�B�@����u�z�\4�ϫ�l��D�3�Q�X
��,��N����Ի�����K�t�\�>���wP�^
>�~�evrs�UBR�D��	��FX�S�h��(ǡ�O�t5殎Etr)�"v�5d9ӡ<E�6z�sqa����N"[�u �~�B_�#�]��y�P4�{���ZO��$�[�c�k��A�M�������>_R������ �8uF�W�1�Ă�F��L�~Ǉ�ю�$�`ʏ�2��hRj�o���@��?l�/}�|D+g49�R�����_^�>�R��V,�y��sE��7QjH���z�����N�i�ܘU�	�3�&24O^=��,�����`ϗɺ�)�p2�c]� �'*w��+d�T
�Fl�EF�����F���Z]I6�'���K�Ա���D�]v	�l�q��=��zN�t�?%'i�&^�.bKk+P�&AtPʼVN%�nב;l��gp�s y`�"��S^��Qv5�M�ŭlhZ��'��D�ç\��qo�T�Ҭ��#x�<o�&�1���>��:|����Xym�(�-y�@�{;C������~j`��^��2>h�?-�=T��~%l����'�M`8�͞�4櫯�� �x��G4 �a/�	���|u�ǗP%�����%.)�59NtO&��H�ՉgiRl�j�gl��u�8�|t&u�I/V�G�5�%@�&8^���)Z`�O��N���-�]�Ŏ=�~wA��g��n�3�Bm����لa�,<sS�w��1�.�ym��FЕF��^�.�h+D��]ԩ�S�L��m�`�)�"5�����(q_�I~��7�  x�ڽz��]A���јqȜ��M^ߍ��m���4�0D�x�T��</c,��)fiɨ�%��??<e-�)�;k;~F;1شXIǾ��S���'�R��B����y.l��W�5 ѱ4�����^�	%�B)�]�Pt�X6�����[�]`�[ v+|��9=�g�P�s�iU��@{�ֱ:c�LTÂ��7�W��^���Od� 5y�ѲpS�'����,)�V4�k5>`sM��|k�,��FO�ɳoo����6_��c�כ�q� �^߇p#[U˷�8�i>Mq@�� �
:|�(�:1B !�o9] K�Ō�F����t6flS�@\�H��[�D��Z*����@�3B�h����a҃�����5OП�:\Ἄ�n�3�'{6��8m�����o��%��J����MU��a���\�U��w-�� ��U�?B���t��	��Pv��0�C�k��P����+(��gn��9\#B�*%�ν�4̽%̪�0�v7=�t����t�W��01�Cg���9�ZG��h�V�r��#�7gh"�x���pc:���)Ä��
���n��)0!]c�&�y�GX	��T�q��%��
����$T�^L��/r#�Hx�W*�5}�(��t]������q�`���9�1�n8�E�=�V;1I�Q� i��A��B�w���U*mN��(�X7�c�@X'�ω�1�����ҭi5���=|�h02 �h��8�5�(�Jj�6��T�S�6�R�I�����l�K-n-�q��ޥ�X���e���&��$�gnԡM�"�f�rsfd�eRKś�Ɋ;�jccхzS��襜��A�wI2���������(�:�۫�I1��y�I,e\]w
��0����������F��<��8~���RD��%��Ϸ�O��.��ң8��D��M���'�u9�f� T5�~��˦��aa�y� ����Ɩ����_.*�ד`�<���}ْ�r�N������8މ���|�,�@|�u�@�����p�
V��SK�a���f��B_�b�X�o�Pp����������w����g���t0�'e8�v���[��0�C�G��u�&�F]�b���OK��q�'X��C��(�gY�DU~�1y�O��=��.��[�6�%}��+��0��`N��P�@�W���j�vF�+a������:�̰�<�����XN�@�*�c���R=�V��5Q�[�%�Q�D�T.�V�&LR�i̞6�=�4��L���7�'�@��OaK1��s���茓��#�M�Ǜ�3u��7�U�(�i׊$���Dcs!�UF���H"�T��a'$2�s��'�-��|}�DH�s���!>R�&V*�g(�w�2�=�HsRkb�4������D�+AF�/d�F��lӍ,W��ڒ;H^z��#��N��W-��Wu�"a�N~s��|���5���5J$�+s�Z�������W-���h|R�yQ}P�p�%��\d���Gc�,��1q�=�0�����<�#���4�W.;(ӜѓXg��nZ�On�F�-(�����TM��G�wC�ɓţ�6#��k(<53wk�s.�vM5�.~�ߣ��!&�-Ac�8]$�*z���i ҈Ǐ��A�lN��l�{�TK����"���rT��AM���3���p�2�z��q;�+�Tܩ>�D�P�;L�o�<�N� �^ ����!������;�R]g�`���m=h�*1�U-q�Yv�@`��\X5}K�s�/��QU8H4vA[a�� }�iADR����r����?\Է�8T"4o��[�2U��y��4�Q��y?g?�FS�NH�&rut�1��W�`�(����!R����$Y���B/�zd��6,��"�*���d�U(p�����=�}�;��Y�@��w�N�I9���sO���;��)��"<<�o���k����.�X��`�e���]��l�ű�;��C!!w@��u���9��_�E)_nR�N^r�=->&l�����	�n
��#�5�A��X�w�����D'�!��"2�� �SS$t/��܆X�a��ӧҜ���b^c��G��v��#(b��d������
��֟��=���I�>��$��X՚p�^p�DG����.�{���`���
�t�/2��j�K�JNPP�n��368r$C�R���R[n;ლ��h��g���� &��Q�6Bඬ��]�h|��$z��d��+.7,Tx��d:�O j�I��ˈL�O�rk5G����=h���� ��vQYi=�nt�ٖa�sp-��[.B~)9hΦ��&����;�n��(�� �*�1��Ϊ����X6�`������o.�1o��Z!YЍ��߲n��)��D�*R:	���]�&4�r�vf�������A(r��d��z6�vMS2����x��#�<���.?�B�oևT�odh9Dr�ۘ��@���h���MJ63�$/ŚU���d���D�*�|���&�!i��d]��W�S͙	�o�FU�Pש$���C��A��,�������q�h�r`!C�̞ljt��{������ȄZ�4��{wc���lq����I�ǌ�x�7��Rm5��~.�7׎Ym(��L^�P$m���}�8;9�<�]-����N3�/�Ԍ�s+w��bz���޵���D�4l�|g=��mi��n�MO�.v�@^��H�T�ᴉ����K���ރ��*#�.�F� �����4�h��� ._.�˭@/�R�F�V������p�a�M���ף���A����bB�W濝酕��R�a�u=��wE4�h�9��2��t)���9,��m�f��ܤ�\�҆���7��Rf���@s_�_� ��gd�(��+���g+�Y���G_g�w�M�^��j��Zۍ&� 7T�g#r���/���0=X��9�.�2��4
N��)�I���^\�J�U��]ǼM�Ջ�ߘ@˵�[*���k������C/Ȅ"v��Ω�OY �(B!E�;sJB�����s���l^8��<�+��ni5&Eh, ;�LΟ_������G.���C��_"�Y�F��*�LO�l�X�[�V�BD8� �K��H��1������o��gu&{(�v��$�Ct��,�NrV�i���}��ToB��`��	(oˬ.FݝU7T��9�<Xˊ��97_���,��}2�=O������ҍ��-��dˬ��t~�nbL[zѺ�5��g��+S��5���bκz���;5@
aG�g�(O�zN�V����W�"������J �O�"�"��5��L
f�h�HM�r��������%	��R!M���#�*�D<� k�� ��]��U$���~Tb����m��7������J�ܲ;7P��q� l����׳(�vu���vw�t�5֭	�Jb*%����4+E�;c��`8j��g6�G��B4SA�y�G��jB�I�<5��h +���F��"P�h�`�N���t�$s �|�W��f� ���?�T�4"�n�Fs��U~>���/��a�!�K`�</75�s�j���0�a�ֵ+)���V��ū�S��fu�#)����rw�F��޾$D�Gw��(��S�\&�u.CN �)��	��T�Ҫ�~�)E�D����84&U�4h)�����F������*a�C���z�<�NM ���S,��hd�@S/'���xwF,𒻪��Ɩ�(���P.�����`,�p�R����+��M�&{yHSk��B ���g�}Ҧb��Db���z#��t��i��;'�+&O��1[6Q-M����
MY�2-�̹�`�]�)�\6!?����,9,�5�C�"�*S�ͫ�N��;�M� O����P���sF�j�+�����G�`h�8�����=��+O�#��t���/Qbd���B|�ŷ[��בHKh�Qh�Vi!AZ�Ps�Wqv�f�	bR�1s�=5�������w
ג���u�L���Zz,�=��tt(�B��!��uP�%O�cHI��� �5F��� ���g�CB�,�o�=�v�e����!}?F*�<��'���ݿ�+՜<m.M���2�B2*m jw�Ƃ���>��/r +�w��iR��2�3�g��Gꌹ���V+������"tN<(��w͇�J���W�|~��֌�2h��p D�^�˴[�� c0�d�+�c����H@�p���z|�"�&���4a�!&Mq��	o���E�Ta�@���u'[��2��T�,��KrE/�ඕ����l��,������MV����Q�!��˔d��D�@�*��v�>=�d��_��ʲY���	�-�U�Ϳ�I�'=  ����3�<��I�ʌ�vUfG+:����S�-$-�.l�(W�H��Ω������O����"��r:�7�7��Q�E�[op�����F��k�cҫ=|졜B�ڳ�M��I���F2OJ���,�$]6܇�
�y���Q}�Z5̜4�b6�O�?�߅<�nR��rͶ�����,������/��'w+�a�P��o��i<�G����?�%���I̡X��pH�;U{�8(�)aC��Ch������s" ��c~%l�c�	�`��$�!�+�&�ofX0MN��l�d� D0.�ܫ��GL���BG��q�?)q]�mǺDvӤ�r�e��󻞇o=q��q2q���5�VW}+�9>is� �\wG*�Y16�j�.1�����Ũ/��_�Y&��{��=�P�/{I����d���pK#�Z���F��c~��=���e�8l���@�Dd��2�>�Ȍ�u�ĳ�ޔ^�GkRS�� x��aG��5�8<��*xco`*�I���]	���V��d��,�qZ:�F���XƽHS&KOg�����hh'�MGG����Q*�;�������,��i��3����s��8�doq�5����T�3i��D�aMtf��=���j�~���Q�����#�:Yk�8�?(���0Y.$�����1�Zәh����B���O��A!��mCw�ٲ@C�יj���c=��z�9��j��"Y\�����[�ð󴝹H�#���������(1te��4ne����i����/�\U&����J��8�SH~�ǫ{i	���+ӣb��J��t�j�p:b6��~��v���Ym�>m��]�����3?��td�nY�����j�wPeLf `	=i�b�V'�[�h�g����t|��C>&�B�4�2��4w��I&R��"�/��x�@�4��U]-�Q���Q�`�>BbK�'�B���I}��V�3Vօz�x#>�i�p�f�thSw��Jb^��� �����$�`��$�E3��m�ʒk󏐼�,�3'g>ح~�66�^<3`�W��i�gayk��b:c��&3<Mf胘���f�(W���ظ��|>�����e�sT�O���������f^&��ڂ5�%Ey
���,�M�>���H��/�p���X���*��ev�a�ģ�2�H��%��T>}�9E�A>���ޭr�(��X.����6� +�wNG%>�I�obv�~4<�����dL�{` !�:@Йq3���~o�6�����2�����8\L�Nf��@�!�N%1,c.��Ed���&��(k	 �D�d|+��TL�m��i��>,�;�}ja�*'�q��k�QI蹍��)A��~������h��{��X���ȿT�,Me:���ե�:���2+�frٿ���U���ޗ�*q'VcO�����+Ⱦ����o2̋�Wz3w�"���KT{x����s�(߄��`�W��zh*y/A��	��xc�\���tZ}��Mv^�Aw)��S"����s�����숯�O��3��rW�~+o��jaԏ�.�80��k0�u�i�<�1p����I���۝�حXR��:F�5o��G�ߚ������OY�Ut�=�d�^ml�ƒ+�+�d��6�����oX�R5
DH��T��K��
��V��B㔉B֊`J�X�NP�?�
��9�2=�'��R�����
�S�{7�cP�5S��bM�v�~G�40꩓�Iǭ6��������N�K^;�xy�9�l��t�:�A���5�M���Ԇ)���i�'n�$�Fo���=ߖ�	W����S0M�M�V����v�Iv���[���6�Py����s����rs>���x�]GV+�v�/Y���D*��C��M��s?⪷@�V�U�׼��k2���:a=p�QA�y�.�FH/~�vxb�)�Q�IX�Hpђ�/�<��;�z��#��3����<�u0�X x@;�؃����$�UU+�1��?�)��+�:��>o�-̬�����TN���[H�<d�P��Ƀl+!P�)�\��Q{ �ӑ�N=sbv��+/~aJ�̊�ߴAgn�b��)jm-�<��|� ƘY^t�%�f~�
i��ݳ�c���0�<m�r8ၱ�Bg#�W��i'��eή�p�kL�ye �#HPho��5$ݎ|
2��X G~q���K�b����D�I����CJ����m:6X
���5f4(4��!�9/_![�=\��O$�u� s�=��$�p�C�2���	wy9S�f$s�ؒP����I�rD�/��@.�M�o��@�~�����ٟ���@)2u��i������V�j'����[����4+�������W��)]=n���xnl7��7�9����g�`�@�y��!;6+�� )n8���9`GG��.��nw����U,_��
�5�x�j������]�8o7_H��.�V�E�n��wu�`5���[�b4�`H^����Jw&���zT���>��+3�Т�\ A�n	zڭ��v'c��Ho����A��4Nxs��(���-^�7B�YF��F���`��l�EL�ʫh�޺�}I���Ow<�E�N���I��ô:'��9�r�*��k�++f��IH�
�̻ȸ����צ"���+{bu;r��0��]0���C۬����F�^z�¿0��7���ٖ<֗���ǹ�N��L����C��*��������C�rW��3����T����EP?����/����:p��g��{S!�L�l�^�F�~�O���͸?�g�t�<"�T������֙��U���&Lp��y�	Z�1�V6k�������A�U���f�͜�h^�֊�Rx��?j�U!?�4S�>&:1|B������U��s��q�v+r$~H����Sl���mr�F� �XHƇa!m�M���uΌ�e��Պ�o�x6�)oK�7:j�ϋM���k���0fI�U�O�BFÄ�^��e?z��Ia������$Y�Кg.����!_\S-���mj�ϲ��n�Ρ��q�v��*B\D��J��Կ'30��(��))���B������Na�q(Ʊ�r[�y��GV��VMR�(�`pS��v#�#c�w�X9��	d��t?�֎�z�Az+��Æ���6���6���U��������a�e-=	�]���=0�e�Q�`�$�]s��u:��|��+�q��J?���k��L��P��ӿ;´�4�;u���h�D�ū��'=�M��-�����oT��l&� 3(iƵ���{�P��/������DRl���*3���qx�CA�V�|J4Ng|�5�����W���k���e�*=;GдM>���>�`��/+��ָ^~e����ԴRV��8>�|�c�:���B��,p(!�F��.a<Y|9G�Sn([Dh�i}O@���(����욬�?Sdդ3�{;l]iî��~�4��Й���A��2���j���0�`���p�&b��օ�Bֽ���_3��]2�\.TOq��a=��`x"/�"\���$�?�c�Б�@��HBI��Lf����*��D�H�}�L%����Ane���G��~�V�1���z���9&Ft��6��p
��@4K��dNT�õhLy����5Sֿ�3��h���_X}+x�Z�O�y|�S-sC����2d���q��'�T�Rvà��C0˵�o��roFd�Pj�	�GH���L��옧A����QT�G�iX�G�w�Wpc�%�okD7E�&�H�K�N�j�����������p��Ǎ�'p�a8��|:Q��+Wtk�����}ثmŦ���v7�C�*Q�!q �oҲGT�e6a�س7f镆��Q��d��U�����z��ٍ��X����[L���j]�"��Q(�6�h�O�
�Pf��0\�e��NO��aB�7���^8�;�H�7Tѽ������Lk�V��ʐ�ƭ���:��D�5X�%�[M��ݑ�Z��ł!�L���n���T2��H�n�x�:���β]X��!�	�xXn"����l�$�cyjqʕWU;�S�`2�|i /���C�O���!I��J]݈���Z��xJ��|U�&׃����h���8���Jo�pr4��<wZ��n��Ah� Uh�g�8��ƀ�x[����Й.x[+@�8��|��i�Ȝ���MŹ��0'��B�hI2�Px�Gi�Ȣ�=���9·X�h)T�w�R�p�b�a0�w���9�?�Л���Cv]V0Qؼ��G����%��p��"���@�*,F{���~/��R�����n��S�Z��s���6��`д�u6U&h�A8�(������?ص�jVM*��G6�p�¢��\A�M�z ���
�LE�Z׸���( n���>J(pd
&�2�K1��"���������	�ݤb����P$�� �oRh|�H��d��`��9�[�&>�#w�f�:��������f#���US���ɎfRZ�n��m�����2��i�g�k�GP�:9<�N�c�|(�=��g��l�<�f��H0E�4�G��b"��l�_G�62I��`L�1*t<nt�rDp�K�e�e���>�I���*X�M��oN�L,��P�v��׵���X��h����qb�B$ʼ��b6�E`�������T����j,"_�o��q�r8�<�D
��3<W�����QJtp�� ����P�d�X4k�nx�܏�H�~b��5p[�>�6�X���>�#_��@����rN�R�V(�Mq����H�	�����DeTX����
N0�i,*�V,ka!n�{y��jj�݆@97<!��H.�Ǫ����:[2Z=���U�X�3널��a 웡[漢8'����7��}�Y������3���$ �<d�$���6a�=ys�zB|:PiӪ�����k�#9M�'�ֆ�	=g�p��F ����O[ۚ.d����
�J�d����n�1�qQZI�0��,i�RE⺜p�(�7wh���%��6�?�5���L�Ǭ�E���P����EP����;��k�@^�-��Ґ�ɕMںF��W��c���<�E��� p7S��$��\�_�c�F�"�F�i?U��H�������T�q�G�k'����yTi�a�銭8�gx������M_�V14�If�i����b�yur]��]��c!�b�-DM�\ȅ?���F����N���
/,��B9�Db����D�T��pGu������9�b�Q�AV_
-�H�(a��Y������U#��8�oQ��8Gz�V(��Zy��^w�-�(<T�)W��Θ{(���l�%Ӡ���nX������i�]�H�̄4d�WB����4{<���I��|�ЂQ����!�&����Z��c7.���5{`}�[��C֠05ZaM���f���>ї��Q,)�V� `�XhNo�_ߖFo��3�}�����w��~��"�ֽ~��Ճe�*[f���Eי��ԧ�8�z">L�MFH�*�>�Ò� g`��;)Q�ίh��~��J�t7�3���U����Y�X ���LɱgbR��p���rqu�jZۉ�y���s�N��;����	F��I-�����t5�� v/��Ȕ��8�Y �'����d���E���Z�h��ђ?�-�uz�t�����C�&�����c灹�����dhP%�H%'!9�@4c�{��s~e���9����!t˄l�p���}�����{/j�-NG�l\��Ro��V�x:��x$x�'��*oLD���:�&�}F�V[+��	L��Ǩ/(����NAk=D��Me/�z �+�����1��$�A������zK4?0�g0Q�č7���g�H�\�?��V)�;��j�!S(Ff�7׸/N��嫈�x#�*��p�n��c*�TzE��P���!G�X/�A��Ɏ_ô�H�&]i_�ݖ��\�$|m}�X��ُ�s&�8��:JV�Ѝu�������z�k�v�X٢�������a
{yDs��0 z�FSX0*���і�����H�hɕ����f���6Q�$!$�OH8�y��m�r�zA��XN^���e�ZnT��������̒2�/�AL����b2�A��9	���H͹nl5��۵D�:y"��U#~|W�۝���e����Eق�`��Y�h��
�6���hiА�q�s�d��Z�е����M����B�}����֧����DD�ґV��y@��*�ؔ���!�)�fD�2��x��%RT�q����tb���>�����c57���lȈPD'
�}�'֛%Ag���o��V��$8��n�O�j���Gгn�֠;.��-pe���AO�r^4��3�"����b����,���q�+��2~� �'.��f53(�?K�o�q��Z�d���2ZGw|n<���7q�u������s�	�i�"�u~lց�pY�Qq+Y�#���#u+[���Q��-(�o5���B�W�Ƞ�ሀ��=��
3x.u&�WQ�I�m���&�̳�a/}�B�o�K������݋}���pzD}�
|e��!�ks\�ͮ��L��O�g�{����w蠉���"v�2KG���==���qT�F���딬9�ה�����M2�j���}�z��D���P���,�h��=�޷^���a�da#z�a:����a8�r�I��m��c�N�]_Q�����`��-��p�0����� �&^�3��.�u6-�u�����u��h��gglXKa�d�DTO����m����{�e�=�i �.����M��¯n0�{!� e��.�_li����~\����������ِk���������I��Ē��G�eF]1=s4�|����{U���ю*�d���IS#[�>����)�h¾ϥ9�?�gT�N9K��>�V��N�cIE�8C�?��i��S����&<UE�O�$-�"�.�գ&Hlz7>Z��6���C���W	�6}�(���K3y�!3���>s� �1c�����"~�qm��.\��/�L^Q�J�%���Tɉ�H���]��u)	P��i���?�D�����HOz�5h��~6�{v��}�VNĝ��j� 0)�#�!��x���L�`�?����(Ψ�-X�}�K�n]����y#z*h���R/E����>�/��3bsT��-_0�H*Tg�����1@�������"ff<2�m��z�Q�P�������΀Jo��h<94q��k�bӥ��
"I�M���f�KW����l�3̧����N���)Av�p�a	���2���E����ހ*�ۖ���T�{��΁�T0������9�
㑨��Jǧ��tڗ�<M�<���sԩT��-���~��#�й%����;p�i�ϼ`�� ��S�J�g]�e�N(Gi�mD�۩w0^�|΁xd	�qw�{��}�O�p~/��v�ƌԦ?�0F��3f�	&�0�HӬ�����ɍ�Y�Ypb��ƭ�vL�	g�L������cn1& �Q����z���xs����!�A�I6���U��ӝ&�]E3n�%"!R(�5Qڪ$"׀|�	�/�܆�\�����x���R�Ͳ� �F����!��7��\&,�k�T���q�.���J�qE��y���~�p'�,��V�r��ŴAQXh�&�s�Uqf8�WYE��x��9�?�R���`��4�v���|�����u�˖�zƼ��!	K㨏�0�#�#vNBP�l�܅HLf��}�D2��j��:�n����:�M6��$�����(�{��,a��j`r�J��j��Z�/�pYm�/�	mڞ��|;��\��l}�]�K�%BO�y�鈿TY`��^�j|a�dN���l���d�DhKH�s�\kl�!�m]��c�۪���'k=3�g8����{L��X&i�a~ ��:;ʑnpw��0�v9�V���>}�r��)�$T^�o��I�`�aL��0�As�:'�P�,����E�:�������ea�D�U�(�~�`�j�.dުp�p��	R�&}!�	QY��x��z�$�;b]���Q-[��P��tߥ�^�߄d]�ք}�sPd!��	����N�|�����y2�ښ*��A�6��o`~�&YE��T��;��u�y�F�d�OP�u�͙G�Wu�ͼ���j��r:�I���nQ"����F �W�~�ɂ(���i���uɖ��\�a����>�����7ZkA�.ɞ�t��z��Y��g�����v�;iR>��"��|�X��gS���}dm�Paء��s?��f�`�N֡� Nq�"1um����\l%���UN�:D��N��+}���W��nQ#��8�E=1��@��Bn.� Ml�uҧ�C&JøCv�Ca���H5�>7mh���g�B���3
P�m#�g�_��s-I�8��\�,Ay�.���?�ʝ/\�@���8��H���~B�	�R���\`_��V�}�����`^ӳ�,�
�+��f�y5�ꕈ��0 ��S��K�o&���=i�< ���X� 3"��КOJV@�Q)f��q��|#�L������S�1���������L��O����sp���?�iQEq΍�-,�+�ɨ�_/���cM�_��\�HO�lӠ���p��T���y`̂��s�� �<�O�e���< ��n��6Z^�̡h�Z��s"g=3�C���g���r��ep�X;9%c�%��?4Na��&�H����Ɂ�~���P���D��ؽ\(P�y_Ύ�2G��n����&쌁�~�)v����t������m��="�r�_���
� �M�q�V���F����Jހ/�@9$��4�b(C A��}ԑl z��_��qӚ�>=�D����X�@,����.6��D�!0/�*�ݬy��
���Ơ5�-Q��LLE�G�Ia�<�j,�[U��>���w��E�F3�\\��T^���a�o�cUw�i$fT��=�)����G_��T%)�+��mc̴�*S��ɵʸߋ�q�w�ƕc��p���(5�>Z�ʍGU��i��5j=����3	I�W3��!�[���7/
_E;�&���:��j��J��<����A�Z�� ���h����UzI LTĽ�V�T�8����7�T��>.�3��@D7+��W̊#?�IN��,V���3���ֶ�0������J��x��#�����jI�We����PM�+�}m��r��Jb�W�F&i��LMs׺"��� ���GQ�|��W`������E��5�]/��hI;Fl��
-�m0Vיk���/��G��U�����<C2̺ȝ���%��kC/	�������<�הu/���R�{�QK��VB�jL�'�}B�)?o�_��J��� @~HbZ���Gf�=U��# ,Y:7����	�s���v�yĹ#Hk�ŋ�k*�s	R?%�T�'�<ǻ<K%��ΉG�Q*I��KPD:��6
�}^SG����*�����(��������6ߞ:��΁�?�N�=#Vmmi0����
�ԛ�+ ����?�?ۜ&|I�W�pBþ�[�(�;����qbu#/��848�2>6Xr���<,���ݡs��v��6���(n[�!���?OB�j�<�t�!��J���r=+����R<�>G16p�������#q����8L���$�G�OV̴�N,r����+ f�Fy�Y��3;�a�[�߃q(�P�I�dl`ӕqN]�5���O%���J#����X�q����?ԍ�B��&�1��<ťj����Z�0R�a�B�ƪ++ʴ��*�|c���:Cl�x�	-Y�3�c����'���31�t+Ӊ�
S�ebb�?�&1l΄	X0`3gB����f�&ԓg������N���nW���Dҳ��nH�,�~4�>W��E_6^��Ʊ�2�?��kR����xHav��� `��þ;�\���n�!����]/���P	7Ǡd���T���m�ꖑ�0s�Z5����}ۇ�}T�tg��R���v�Wrҟ`�o��aS�k��;�%ey���KUl�hy�e���V��w"Ln���q�o*)-~gj�ri�V��w-ѽ� �&����<��ؗ炥�o"��2�T)���t�6}e�x��̮j��wg�r���������!_n_$�6R���cU3t�;�(gzj��W�w7Ag��R�Z�~s*j�W�۴�'�t���hRĘ���<ř�AE�S����%�&[�f��!AW ��t`"�:���[�Z�hy.!??l\�Cȳ	7��|���1u��\����5KG�J��l��.�-SfG�#u�T9_% ?�Fn?�4LN�"���9��P�𝯇P �Gp���|�<�g���N�'�Ф\?�Ar��(�7��b]bMmrR�W`�Oc<�����{�PvH���bƱ �����m��Y= ���P��B�q��*�i	f��i�V �v���AYѭ�w)Az2s���	��H���9'�N�'�)�)!ݨ�!џPT��L��Z	(+
���ߎ�(��0ꎝ� 2�����sX�A,*2pӂ�uW$�rU!�	t���_s8�=(qX*�|*�{��jZ�B��k޾9D��=o���
�s��p#6�S�pAD^�R�V�����_�A��߄�P,a��?<zW�a�;�l�����p�I���f��=>D�WUR�$��k�C�`�xp�u�(��=����b�k��/m!Pgy�Ifj;�`<�g���Bxp��o��$3�İ�jU��C�o*Hs<*���
��V���_��H�X��\��AÕwq��K��s��T�	�\w���55$8]��C���C~�@t0}��/W��y�[�r!Ӂ�˔��2�?�I�v &T �p|���1�j��`pd�?5�B�><M��9~���	�v��դqo�ˣ�m��f�Y޶������-+�S5�1+̯�^+i`P� �P���U��k��v�<�.&ן.7�,dg�H��.����.����#{�S���ƐX�i��@u�
���h�ˬѮ���X���5 �[��ϣ�
B�\갦�+��+ gA�l>Ϟ�%`Rε�~w����m�9V�J����Ԇ����ѵ$- �8� ���P���m�0'���Β�u[�e�cɬʘ��E�yrՉ�j(+Rz*��΂�^a 4x�i�i	� G,�M���>�/Ebh��S� �{O{@�jw#�h�UpL�����h��4�R6^>�ܚ����I�Je=N���{<�E����H�,gB I9Z]�m6�͛c�9���;��>K=�+cL^U�����/�Tw�6�ɛ�g����M��bSW�HYi �\�qf��z��kb�O� �L����u��4o��Ͳ�[������{0�����^�?�9����-9k�����^#�m0ш��s{�x�^�»+�_Q]Nb��#�
$��y��+gɠ	��!�e'k����=LT<]�O>1p^�<e�{
� �Z%��YT��90���� ��ha�0��������+F��a����"Gcz߶�O� �q���vKP �������]�(��ڤ3��ȵ�D�$t$�h؊Q�Zݢ�L��Q�{����P���#�1����=�]���w�l������C�u5!%�����,�_��:�7^�>l٩�\����n����'���s��M���N���;�,*�@4��v�A�7/�t쎻?���=�=>ט�׃��y���@5��Z�q��2�.�̽p�:k�*��0�Z����vo�$�~�~U�v�d���i��J9����/��z�5���kl`D�f�Ȍ$��t�Fg��v :a�*��>��b��]�x��ޥ�TD!��,�M�4lg��'߲#�9�Ӿ��qF%Q�I�O�1=cj��<�]��s���� �P��%n�{`�%(MP:�z���,�^:7�q2�g��-_�1��i�qIl���gYR!(�V��$��o�~!t*=��2D�S;0=A�3��w�a�g�E2�[��Ԍ9%W��V���+k�r@o1�Œi�.���1��(�u��l�v�e<pPL�̵�)4��GȫX▟������(�e��v����<'+�6���~E��\�������4������+ �3H��I�x�`�bdТ�^ݞkV�2:�<�>,�c� 9�Ȯ������р�)�78^�Q�\%WV:L�{�tq}��v�6E�X�*���_��:܂�-�Tvk��+|tp.�ɺ0t{`��7Vt����(R�$0�'�J%��Ǒ�Z�U�sn���v8�,m��D�y�!3�.;��A�%t�eG�6Tr���+j���[2@�6tx�1�$���k׋�Z�Q��5�I��w�s�M&�p��=+�r�yT�h����䖽�#fY5�`i2Eu��wV#_��w�����'s9J:�VC��)�
�����A:+���e��t�_��N*��B���T_��<c�,;�^�>H�?EȅQ��9)I��鶼����4�.�	�h^ѷ�U�Ĵ��Q��� �z��t�+ۋ��oV��؜���SP&.�)#8 2�Ǘ�\*&��x%bg�d�)?7	R@����Ĵ����L1J|i{�H󭇛�9�;@��nV|��T2�f5a�m��2��G(Z����֡�q�����Ѳ�dc.�;+>;9�_d���JN�貆T�aR�\h��F@�˷������V�շX�ƿ��W��V�9�"�[:��|Ǘ}����/O�b�9�Tg��4- .c�W������/�/>�%C���Me��E;����ط���+y�!��d����YA���qv,kó��'������Q�Q��W�?� u�o��F�9A�R���\���2����z�h���1�X��W��J���۳N ��� ��P�8v����)@i ��q8hG��@�k� �BytQ,� ;~F~���Y�w����>9 ASB��<*���8�7�ǫ���S��G�'$���K����M�z�>��1���ٷRx?{���ν"w��T;�#+��o�[���މ�н3�٘����!�vO닪�������a���4�5h�k��̯8���0;�G�~��IA�|D�co�: ��_;�z{�1&����]�4��]`#�j���a_�>~c\BJ�#�ϳ{�/p�$�}pG^��"G^�*PB
3�0a��S2+ٞ��'=�\��d� s>��_3P�����0�����A:���S٧�V���K���!��֣�xP��UҼ��A� O�#,�$j���{J_�L$�68?'m��'�Ǿ��͌ճ�G�9r�*t-	��;���
�c*�I��PG���ƈ�Q���>���P�A6�ѱ��o!�(hg��ٞAWx�GW�l����
���?wo����e	�Q������W_�?��I�d'�.@�%[m6'�U�$ǔ+�nUL���5��>�MF���E���1�~x2A]#7ꂎ?r"7Z,�i�5��nk�����x���r,�{�v9��'B,���W���1�����������۵<s*G�v�x�J�n��*����k1�(�	�f���͕��=������y����n'C����yk'�֎�f�����{_�g��! ���9&��#��'�17rͬ�!�������sC��w�����wToX�e=cL��/�J�Lݟ�r�<\=+߿�0p�)ś�䳘 ۨ���D���U�x0����ԇ��_N��c�1�p�}:%�*��#p���z��4�{�5�'�#vⶎ�r��ۈ��x&u��dO�_2fA�+C�3͝�T$��!�.�`���D��x��4�B�ٚ���..�e@���e5�D��=�ޖ�3eT���"���/�B�)������n���� )���a��FH�bzF|�8@ճ%f��3{ ��[��k���2ݤ���)S���}�Kw G@d���e4`����ݵ�h��b@u�vJ�;���@0����"R�čB�>����j%�$���%5=)Fƅ,6M�g�*��pc�~���Ӂ�jC�K���,���}�XQ`¾���;����� �̒Ht8#�/I,�L��3~5��E�L������2��t����oz8iL��Q�ި]��v}!��a^M��u%�����zK}l���'&�fB�+GL���e����f���M2�L�u{���z���K,TLm%��V\�Jc��	ؔ���^x	z3�C�v�S.[��ms��{�/�zZ�����:�Ɋ��cI޽�����S�* cWԮ4���F�T�dv�j~�R^}����:���'݇�7TP�u ��G�C���H_S���V n��M�}|�i"Cl�K@��hа�I�%�=�z�=�U'MI�qI1�6�����P�,M=L�S��mFAJ�1��lzt���{��3dwN��b	r*  7<��FVe�~���P7����Fx�S����H��?�~��,����S �q�I�����.��"�(_��%Sv�Ώ������b���*����Y�atV/�GY�~�~D��l[�_����5����v��UtF��
�"�g,G��-C譄���ǱO���^�oj�Ё�;kT4����ᝫ_y#��x{�҃�P��dl���AM5Ύg��*O�(m�������y��
n�I?��/^a ��ƷP+ ȉ���$��5hcO�]ӌ]W�HA����Fm��o"�J��O�M�lkˠ*�'�,��h��M�
: �(R���ӯ��6�X�X@�{��w�fWO	16K"r�����v��>X홌.i�#Y*F6��)R�N%�P$�ѱc���־���}��cn�'�_a�q���o�t�`0H �e��_��f"��xF�ƲB�+c���bi�������~<gG�1���Q�WWg=b�}��@B�֖�"�Dy�2��uT����&(�%���%D���ҽ�=�-��[����v��P��>M����,~�����#��A۴)^�w��쎔��qB�E�MeF�<�sra	�ٓ��0�I��cշX��Or�nQ�-�M�z�D����/�blꚠ�E>���u�O-�3��+Tn�{u�~�drESy������i�0�&eléM`����.�D��ve֨a���EimM�ܯe��4Vv�]@����+m4L�Ӂ���P��Rݰ��7����]]�F3
Ĵ
���M�͘��9@��ЭAI:g�� �~V-}�_f������1��Y3��G(���1�|����&���G-`Dt�)��2IE����-�k�E=`k����Sӣ~��K��g�w�x��P�H���g�e����>�����zQJ����-�4��&�t�y8�xXg��: *�k��5�9���"Gj����j�ѵ��=n�P,4*-LI�}1�X΍�	���r���i��C%�6\F\QQ���7v�m31>�v�����fI��\��:'a|&�뱡�*���E�j����ɡ1���=��S�� ��j�;�}816�8E�z�x6�$�ʻ�ߘzc��[3<��k���� �=e�F%Jp7�K��V���j��U ���C�Y�FR�����soO\'/��1�p���Mbm�'u�h�ʁɁ�Qoh���r�P7h􂦲@[�/EC�?�y�9�2������r-�C���<�#�-�>{�Wi�*����͓�XDb:�8�hl8���B���9I�F��|�R��ʕuy螥� |�!���i$�]���B�L7��l��F]X�� �Uے[,b���ܬ̑죌���f�Z�y�Ʀ��) ��_h�*CG&�:�{x��>�g(����d�!!�W��� �,�P~�/�c�/�{�5�-|/aL�@:b�$��o��.3 ��o�fd��Zm���]VF��Cn�9��j�JC�>�4U������ G'�	��yc"��T�O[W��I8�\� 	T���=C��$��愪DA�//
�/�h��9���vS����_�_�?Mf����Ì�0����6�Q�V�^��+4�]�1��!���GH�Q�3������
}�`�N�*�4D�W�Df��`��]	�F��|T�D�T�S����J�1

5ɟA-߸�!s!R�:?'ϯ"���6K[oT���o�h�?u"0�m��g�^���3-2��x|FG�,�*s�D��ʀÖ�A�/�s�}���a��h�;��|��4�r��R�(�o�x�Q��))ZD�m�a�I1���(�á�G2�	��G���^F��I�ѐ��{�����=��:ON�Fs��p-[賏��|����tdlM�J�� �Bqm<��Ez{��ǿ�X��3�֑���Qn�g���K2N���U����T���������?�û� ����B�B󷓡$�u����U�<{1cx�����A ��X�Q�szo�m:!n��D�����v�C�<vΰK���QiIT��?�,����׀mc��@����P�QMsL����0 ��^=¨�3�^(@5�(ƚr�ڱ�j3f��Ea %�u���C[�q8�KS|l23���T�Ws|�b$�(���%3��kvN`4T���d�����iA,"�1W��`�>����Ec�	K��J�#/� ���}t��_Z��#�tt�z��ۨ�xCN�a���9#������M$3��v�p|x������ن��k�
ڒ�6a/lA��<r�`�]E?[��8l�Sz�m��B� F:r��R��=��t'GO��_�Ž�xe��rj�=�e�9?<��N���F�'�C�������g|Cn�����>��`?6E���N�J��@�*�59�㤾��Y�����:�"�@q6v;ZuV�Z��0��MS\�Yk�*kI����$�"	ztB�%���N��4飖�U$��wwܥf�k��/��@l�dS��	���ӟ/1ГR��2�VW>(*Pʟ����u�1��9<�sm ^bw0�JX�
�H�6�`:�V[�N��Rs����pw��m�cS��'4
V����T��� r�|�x~����t��^�=�'y	pF�v�=bz[�=�Z͟�gZaj��}��r�%�WhK�$�f"�Y9�U�W�98}�O��;�TB�'޷�"�/�����+�f�©i��Kʳ��N����IO4	j�9�I2�
�FÃ�ᔔ��U�����(��*����5	�H$�'(����Jل�<2�������ppd�{�������5��������+�Y�X5zI���M�x��6u]���[(�F�}1���S��Id�z�uV�4��&
�i����K^g.qܬ]x���ȝ�h��f86��T�� �-4��c��l�����i�ҙjM���ՠ���,[yz͝�����\��]���q�"30��&�C[m�6O܍��7
J��nEV��q�e,��V�9}o&Q�į%U8�X7��0y�T�(@�\����A�7$ϐ�T]� 03c�'Σ���C�{��d�n2ҷ���y<��!��_	Q0���l#T��;�D}͆�y��*L<���f?�ǹ5AQ����6�����f��i��[0��&�lF�3��J{�=)�6/�0N9�+x'�=)���>c�Ȼ����GaÐ�9�<��~��@��`����@��A�5o_��W��)�G�^L@F$��J��z��G+���y�3pj��!o�2��nX����ŷ�k2�����d�9��9F��
��a�i\�^$��ه�+�5���*�[D#�J���~'�Ɔ|��Z�p��Y�/3�3�J��L�\������px�����"婅]@fn�#R*A�W�U'q�?��y����C��A�IYP��ю�W<�O/�l	"i�"���&#d96�ɠ.lvI�:Ľؼ~�w�I�gT�_&ț�ح�̙r�����` ���w`56ﮠ�w�h��!��Z��C�O�ob7�K|��%��A�F��@6x`V�,���&�>�m�+�
�};4�Z��f%[MT�6���d���%�J6��z���]Ϯ�+¯~ٷTU�"�P�Y�̗����^-�����i/�=��G��6���x`Kz��yV����鴭�$2�ڐ�K����&��XTF�[5<M&s��k���}"�Q�0u�w"	뗤}H��)�����`�:�P=�K!�i/���T�W',��T%o8�phw]�u�Fp�����z�v�#?fl��߄��i��� ��j<wDf��^ � ��5#9T�p<�;7�FtM pӸ�-����4����b����5�@�tH�8�_B,ߙ3�ySn�������礞��Je �
<߿��d�7��1%fѼN6:cu���$���Rs������_��[1�C/�=�oy����ZXE]_Cǟ@:���غ��o��ǉAY{���M��W�K�PأO� |����k�"svr��u'X�E/[��8"B�HQ��Y;���p�X)}�j�a�@(�P���Ҧ~���7Ԗ�H�o:��W�;��0��IaҼ|�|Nx%._R�gʞ��W�qvNK2c�e/���K	������
i�M�m0� �g��$	Lt�(O�"��������>�<_ � �t��/��tR��z��A7�K�b'ֹ�߼�2S��	H��@�t�j��Gt���E�S�Y��6��	�R$���U�s�X���������_�0y2E|.jh$_ ���f�T�1����!w�X��[����:���͕��!�� ����=1	��f��#{K�Bd	�����8]N�����	��!�K�a'4�Y�\~�K��D�lL>W����d�z���ܕI��#ObD1��e���,i>ijc�Y�k^gd5�:�<���\������ON�Qj�5�W�!��S
l��aT��h��6�'��#�y��U��@�K��@�)Wg�"� $�1��iJ8ׁ���W�eWFÅpo9��[6o��3��!6.��o_����2���GX���oI}���#�mIG$+���t3�O�1��^�l�`Me|T�B�$|�ڞ/�n	 (��v�̙����������R�8��۹�E��؂�_�F����6�ź>�D���:��[2�`N���Xl!bR�R } oc�`�fE%krp�Nvo1A��ߪ�����>zu�G<��uA��C�)/h���t���绺�A5K�r�/c~Lx���
�Q!Y�����D��b������ݦ�5����L����!I�~���s��+n�qj��pqG㔲�\m�����ͧ�I�f���� 0�����v֕>Y2�{T��8�2����w@D��7FE)�g��8�H�Œ����Ct"���K29�9v�u��������ع���JO%��("����d�q��b-T^��̗�������T(l��P�Ƭݫ�v ��t{bo䊏�K�rf�'N<-i<���:B��s��ĕG�W�[�XVы0��g���n̔ᄀύ�h����$��;�c�>�[��G���J����ɷ��N�AbW��5)x�AFks.�d�*&�����և��m�t�!#��Q�g�������<�ocs����8|�D�QkaF�\�+�"Q�-��b��5�#Bl$���$�C�f\�����&������}��*V8c���/�Y��J�P0�My��yR�k��1y;�n��
`읒W%�#��󕦚CH�,t`��;��њ ���1� K�����U�gS"kS�z�=��S,� �e�u��E����~��6�e��f������?���2�]NL�
�K�#��R��tl%��y4g}�%=)�>��;�Z���`샫f6ψW���0�-U�%�"�b4����.��x�4�0$��4j�L��0.a�D�r�exB���J�I��	Z�k�	��s�fT����pG�vb��v���v�)�ly-�[L5�넋�f��z�&b��u�^]'���Q��AI��n0j�9�x4�;�����Z79�1���v�ָ�໱����̅�$��i{���nO?v�d��`NUL����1m�1P�T��0��b�Ъ��2�����@V"�sC|�2���	;�36"+�@Tg̈́��ols��l���짬'�+=��_�1�i����A�N,y^g��n��NN�W����΄4C`&�/:���Ct��(ӟ��Q؃�^��$�dt���@���7��-Vm|N?0���M���1^0��6�c��bD���8H�V)m{دg�Q]���@�d�Y����ʢ��HyL��aX�?֍�Cv[hл��R�����`�gy���A��lf����ml+��^۶�K��Sg�l���]�F�J�9��8�R��.Ţ�����2�ǘ�
Hx� ��Z|B�x�ǆD)�Eđ2B��_��s(#��^3}��Di��6��-��NF��_J��P#�4K/dM�Z�1�h���¹Z�+����;�H<Sk,<w"ߝ��/fԻ�|��8�T��=�#Q�7N{^��2����~���n3�t��G�m�x�W@�ռץ*�_�^�59j�����^%խd��FS�zgs��oOG�"i��R'2�XL��+��N����+H���Y����)ڽRc w�U�\�YD.�?	�K����)��㚻P;nP���v*`q42�?��<�:C����;�ko$�mi{t�!
0/��h���wϷͿ�<B��A�����r��㦚`�4sO�°�-��{*��������xY1�;��J�2��$Q~/|(��_�\��xxAW6}͵Tf6<�vS]�3Ӯ"�J 1��ƭIL�>�����kN�!3�t����������z����s�J�a�HN����d�s�
��
	��"��^:>-�r�����gc��иi1�Z^^Lvd�-^2Hj�VW�֠/�@�	���v@�|�$"�Wڗ
�M����6-�3�{`n��Y9)�h����_���̞��J�Ui��Q���$�5��͇F_:��KϦ ۻ8��zߕ��|�2N&,;N��yv:y�
6p������?�c[�!KfbMO I�Vud��_���
.*�X)�n��ê�;a����k��2ĸ�Le1I��\�	�v��R�Qg~��qLV�b�h�r���t�ЎS��7���I��P���}e�����l���z�#%FH���إI��j�4,����Ã"~<�,ul��ݟ�ڋ`C(K�^�Q�	JU�%���׻xk�T�4B\�W��CG.�_��la�c�K����sY�d`�r��ب�η�9Il�W�A ��L�2Q�-ċ���V��N��|��N����-��5a���$8�\��;����$j���[$u�r�h�}�>�Ne��Y�m�w0�
V�K���� �{��u�\*�aq�"�q55+�^�'��6���b�i�kנ/�*N��b`z9�ĸ2mbEs �<��X�������s�$���;�z�5�t�V�w�~0��!0+}���oF��4Y3�E,Q�#�'�6o]��Xs3����Qca���Y�F���c�|������"��[��՛?lV?��<Wsf\1f�ҎC��N����h9�,
)/������p	�м�W7�j�|S��ͽ}��Y�n)3y*"��'%�KvaϮ���uZ��-}��g��sE
��z<~�soho��Փ���m�6�K��m1���)�Wb{�nF�A=��?����4��H�@V�x�g�Ct��4�� � �f9����#
��0䶃�%�pʽ9}C�B�Lo�B�a�}�u�{ l;�_� =r�!͆k�o�x��j+�v�"a,od x�]�� �\�D�IE��ǰ�.����Bx��&М�31k�p��W����
$DPIa�9>�����{�ᬝ��bb���WB�����$k��b�;G�d#�W����S�,����3��'%}ǌ�^�n8#�!}b�+� ���ۈG#P;::`�����yf�PΆ���F���y�Б�լ4���P�[ǥ��V`qʲ�}��_h���w<r��lb�㰈�_z����X�2�/���8�p61'Y.�����_rmT �&w��E#zVt�S�%�C���eD�:�#-��J�x��⫞6��J��$�X��U�U[�=)���䌱��c[I�t�� =h�{�B��lV�W�����b ��vj���i��P���L4��Ķ=��|�ID�^�9�E[���:o�m�}�y�w/)F5�[���t>
ݛ�n�d`5P��ɝ�zr=y�#̾�QX����뜼�Utጊ<,��_%���x\�ғI�'-eM�bq mmi�)�0/�.�/߭~��4�U'ƭ=A�b��h�ˍ�'�"�Q����U�خ�Rp���DE��TQ�;�*^�]B@"u���2£����ݹ����YJ���� ��~�4O�(:��>p��n���2�~�r<?G҈2�&1k�ST��q����%���Tn`{n���}��X���hTr/�
?�/y�NSY`1#}�U��T/5)
��,6�W���Lb:)gk�~.,��X��_2Q3ǟ�<�/Ui����|��PP��\�RFWI%��S珡��1^+��.{��w=�ͣX�E/�Ʊ��ן�Z6+��:��~e<,
�c�7ߋ~X��i�8�]Dh�L�pzO!�Ǟ3jp��ն�[�7�M*�x4)*��A:8��TųqZ��E��u;qwq��յdE=�s�j���9� ��"�Nu߯��y����]�F!&3��~�-G�d)d�'�t^q���zSP�������J��'�f9��W]�ďX�A��qe�yL���d��%��77>jr����%�[��R��"�q�_����C�����g<#%Kj�Xu��^�X�����_B�h�2p�BTx��ʝ��Ε��'��+���D$��Z�K�Mދ}�}y>��oEH��!�6-;� �����K��-�	skIX�ﳶ�7l܃o�%=B+T�~3�h5��Q��iW�Ҩ�ߴ1	�J���S�,����&	{�,�f�����n��G�*����Q�yv/�a�7�W��g� H�m:�3�G�W+M��&�+��ߐ7+��mj�6 Í�u�G�+X\�t�\g���R�e�h���W04E�YQz�E��_�B5d��J����0� R/W0n��B[�F�}��|�����nԼ�[^��A�'����t%��hD8ݩ��)N�1{
����^U��<c���k�>"��it��P%\#*��� �u��S{�/�-�����n�sJ��Q,X��#\���O0'J}��?�P1b`R���'5r[_ ��ܨW��y����Zs[�$c8��rT��� o�Y	���*HO�uΨ�k)&Ҁa�A�d0X>-�<ռ.�y��q�V��l�zd0���Uo[�y�]���ߡ���9H�%s>*F�rE���������n��؀��C�tɱ���J�\�{0l��YNq��#(@['88�Yx��1��:aiׇ�٢ _#�/���4tGjM«g>��+�G��4�P�6�1n��߀4���km�z�I���g���X]�_�5>��"1�uN���̳�o�P|<Á��׸Z��Xg�2�s�,���a#C��������>R�hw��C"���`X�����&�E�+ Ns
k��K�]��ó��"��֭�.0��͓EZ:�r�G
�6�Ò��ެd�c�W���^FA �S��{�KZ��g�f2�HȦ�nhn��6:r{9_�����Yb�T��&s�0��5EQ�ov1yb�)b���&��F@j�^+�2��cb	UF0x�
����-9�؝��W�'�%��b�t&�����|���l�;ք�ݏ�TyCW3�@��
j��R�ܭ�0L8S�U��Wr9�M,g�b�o)o��"YΑ�j��Q� x��dk�����z�������;�A�P^��֏�x�J1k~�<i+,w|�G�F��8Gg�q�����Q2-������/��{���;Y��o%B���{�����/0��3�&�o�S+V�~���H�$ҍ��\�i���O��"?��oBZ���qtP�L��5�%�G���/���j�����3��Ҁ�{D�k&��Hz�i�GK�B�d	ma�m�'aM��@���F�3X ���.Z���E�,<S�nRg�s��	|�>�J��N�&G�m�����a^*�h9Ƨ�����>cJ>�Wk��Z%C��߆ث�#�u��')�c�PZ�0��c{f�ac��]��?�Nq�����5�}amZ�X�:=�v⬺a��C�x!f�C�a��N���*����(J+a�l��\[pƣ�i�m_O������W���O���M]�N���c{N�(�W*�\�#`�Cp������VK+[���ڊ�{L�\f%�ಯ?����x��~I�1�]��y����Ej����{c�+�d��v�]����6|P��Da1zM�?�;}��)�9��l��G�� ����y��!;
wPٖ��ٽC`��##R�ܰ�<ƆՇ�%1�G��t���6|E���P� M.�ګE5�?P���7�<E��ପ�7!��9h37%}q$c���4�}%%�W�9�<�~U~4��(� �hj����۠ &�` �*e����,l���D���WE��^`[{X�M���f�T(�6���Y��fc�'D5`\iGo-���̿|\��,<�=����x�c��b�e�xA&�ƣ_Mz��]�V����k�mz9��t��znh�|�M�kP���(��Ȅ���`����i��&W#��0�V�g�r�zǻP�s:�h���-��!�
3���S��Xo���4�*ˊ>��2��T�h��?��C�a[����'{���
��s�T`�.q���45�]ݽ�	A�K����Ɯ�Z��o`^��'��ڭ��ȫ���n�Y�'���ƺ-�t�X1L�5�o���'��j��iE�<b1&,-�v	�5��B�@���~����~�L�[��*��H�����xJBI�`b�2���\����II��K������7���\��%�N��~��&
��Z�k��f	�_
�"(��{�JW�c<�ӺLIQwғ*x8@��?�����=ƀH"7�KG��������l����H�?��V_�/�r�+Y��0y( H"�qf�2�b�������p���'vzL��'{�;�Q��E9��^J]����<�eI�����gxz'��\4筊l�y��f��|܋���M�u��k0e��8n�ĭh��I�i0h�
����.��N^b��9!H�u�-H�o�V7(�P}]�q�5Y� _o�.���i��5�Ǿ��P��7�[8����W�+�^��W���瓴��e}����R������X,��T���F��7|q��L�/=p�JӑGx1��%+�z9�X
k�/E���l�&�H��boV"�w���,�JJ ��/w���`Sk�/"B�H;09�ֻὯ�����kSp�k,�up#�u����א�������|�ގ��=�����J�٣�@+�ӟ��q��wS���}�z1�/\��SR+�[y��m\��HPhsj]Y��e�g�z�";�|�ĺɘ��q��� 8��7s��q��ｄ�.R���ރ�ӸP
f������:S�U9��(B���	Ǡ�i}����ה�+] eV-�+��e9�#�6y�1��ql@�#յu�l;��d�&�m�����,�6�َ��+�8t�ŉTiښf���*>	�����(q�i��Q������5M�����¥�QϺp��(�y��&C�=�%~��	�NNh�2��&��s�������V5��'���)Ɲ#�b��K�a��wS]� Sx�z���V��ǛZ�h�
�f�ޡ�	���Yr6V�'�����e1�Q�~���H�=�lF(՝�8��f��-U����x5�5U@{x3�T#�#}i�v���I���Y{{m��?��μ]6Ё��w`dM7�q=e�k��m��pzg_�2�<$�^�>AC��J��6K�{�ս���ß�ٝ��]ӑ�l4y|˾O��G�:0���Ë_�I�B����mJ0�i���^�(x
e�E�Q� �Y4D{��Fw�����1	aZ�e	��}g�Ֆ(m`-��p�-;ƀ}�L񊘋���Ȭ#'J�v7
a�o� ���AH}�^��-Y�Y� �cuZ���*8B���cWK��4"xv�-�ʂS�Q��GW�ً�%}�?&���L�Cc�s�s�0+*����+w�''�F�\��&����-.6�;�V���\��A0h�%p�gN���-�ح�������ۋ�fם\uB��H!t������*vM����F���*npNT�]h�OEw�%
�s�-=�9ﵼF.��0�M.��)�f�Jr�c�����������^"U���l-�6=�,�td�����evM�u��T�)�1���0���Z]:(��XY�Y�0�*��Z��Q�W���xG�	�1�D�G���%a�b��*!�>1�R���f��ρ�W��o�F��+kh���>6A�K���:`�m�/�Y8�z�GWgCb��n=�;�!;��64���I�v�ܵ��s�f�P��?է�ɬ�I]�9QJ�3�{C��Ӕ���9ٰ{�Ȥ���^����\7��^1호�g�^&�����E���RK���:T����D�)�3��VB��e�%��=��͖��Sl ����'�HN$��&+���,�25G�1ް�%�����^ZJ��ӏ�?�	;�lM�Po6\������C�kXf实�a�:[�G�]�DG�u9I��!�^p�O�ҙ��?�S��I>�Κ�C/����렩�T6 �%���������$u�?Jv:����$qe���C^�`vK�j�gMxV�L5�`l�dwzA*�^��b��;�'�;m��d����Xe�4e��a[胤�u�?)�?���S�Xq1UH�Û�-�0��t�ܨ%�Шe����B��w��03���ͭ���f��Q�i�;�rS�r<w��ڙ>�OSL&����?h� V0��IB�w��ҍ��A+��yN��]�;�Ǘ\A�-!��s�Tn�-�}`��[Iz2#�ܴL.w��m���|��/���Iy(u�E�ul^��Z8�[�<}�\�E�g�!.h�½�T]^���Q����O��D|2�P��,��/:f�G���6��0W�h��P7��r�}���AY�=v�}���;OH���1[^���w�������W��۱�S�r<�2i4y�ս���$��Ց��z]c{~��g��ۍ)�i9���g�p�[C��Y���	ە�e3h>�'<r�_���Q��x��z�K�ì�AN�,���ޅdQ����*��[�g�*V�"!�4I��Ģ�����u�0h�o*�U�k���Cb?��lt��S��k�e���v/����Z�:�	������ƥ�8Q�&0i
i��T~d�T!F��NC�RA!]_�LDĝ��K�Bif%L�1ܑ�,~�y��,���o�S�2�X���Ƨ�{�yZ�T�4R!�ɭE|K�(0�z�è�:������!f��-��^�*c��Xވ*�HT���7o�]v�)��I�B�#P|-ҭ�x2mH�`��G��\�`A>����OJ���j{:�t�|��*j](�x�)2!]�^��:���Sg����tN2 QKk� ۘ悀�c"���9	D�:^(�Y��j
A����5�G^��G�6u��^
}�r%
棸(��a3��=������ ˰�,fH7���8D۰ހ)�G�;�Er��1bE�7vN�c��RL�7u�kL���L�ke[M����l�ҍʫZ��'b$c���1���A�)�n�E5�U�\��XD�)u%�!�9�{���Ř/tz`)C���0���G˪��
7�%{�[,\YAVhp�Hۊ|��g���!mN &5�ih�U�[| �h�v�7t�����$��J�r�ۭڝC(ζ��<D�Ǎ2��ǚN� �ixV�yXpQEV�����SvE�0v��Msl�
1a�����"홾���'��Øb�AGe�J$���Ѱ�=�<X��S����*�,���[Z��D^�'�z�:�~8�X0��z WY�nwy`|�3�IX��{�Hs�a_m�!�v�,!�շ@7/
�+g��h� ���H�kl(ɻ��i�g�\W�L�q��G��<E#.u���b�=��[20N�cɆaG�x/pNh�4�w�\�)�-���Nj,�8�}
�+��Z�q�8��@%���S��eSx���ǐ"+�'d�����<zD�1�+/��ψ����p��Ud�Sް-ŀ��2x��+A9 �����6�s(�Y�ޝ�����������:���\@Ű����Yja�D8�
�����wY���~V�V�b,���T4u���H0�vQ3���pı��8�b�硭c[��&�M��7��~��~�Y!�O�}��
�Ia8� �e��-*ϝ��|_��K�D�m�������!�J"����W���4�oD#l�Dkw��/T�u|�67p"����1���d)1����p�ȱ�s��P��+��'f3�D����ϕe�Lߊ[f�I�����H��h	M�D�� � ���2�5�ZSe�� t�7\]�;ӋxV@�,"q�F��O'���*��wp�wm�|l3/��]�-�D(�-�b�� ��$#ξ����|��M�3B%fV�$��牰A��0���O1�i��OD^Ǎ���T�s���g��F�oH��}�8�#��P��Y.hM�T������tܾv`�V1FbEV&��^y\t�t�:~�)W�M9���<v�+����l1X~!�pt��h�:4��t~%�u��8V��}<��˔��C�C�#Jk�,d�y(��o9\yq	t^*3����)ږU�N�A�}�^�pp���Ȝ���W����{~&4;�Y^+���� �.E�� �� �&����o�b�eiC((�Z�e>�<N����&�t��{�G�%��7�ؖML�=Q��.���C�8�5#ZQ$���̯s��v�0R"*�K���T4aӷor����&��F.���qҬS(�Sѐ+�&l6>o�*=Sq��2�9{��D��	DvU᫄�(��#� ��I�b�&4�U��q\]9�@WH޿�H���-!�����7�?�+��B�����X�� �1�ě2sL�ꐔRj뚂6�]�gى��n0��7x`Q^�2����'K���x[�Hq��Z.�uΣ���4AI�ۖd�J��ҟ��N͵8� 6=���P+b{�T��oZܞ���YXx	��#j���Kp��y��ZW�qaWU9���	��#�2�����4��� ���݈�Ei�i�2-������������3��R`�mͲ�j��2��?��UCNcz-��� ȟ�� ��/�F���o��6>cjC�+��8�w�ΈY�u�oa�)qN�8�+�^η�T�
;�����;���ӿ����C-K�i���H���t���m��3� �/J��^}�����|b�L$��H�r1��<H�nz�j=_��!`4v����ث@盧�t�FG�BlTɔ�l�u��ɪ=a�rs&$�x^�#%�RD�犟#�+z2��'Sg0j�c���3���Y��@�����j�8r�o�'�{VgI��C�$��t��x�;�	�U���Y���^��!����X$�.��Ȯ.}�Z���3-Ao�s$k{@��G��Qe����=�t�j�`��(>�Og�7	dt�-�SdZ
��1t��6�|߾�����0Iw���]��H��ԕ�� 0K�����Mц�2���� �"�r��K�DzM�@F�ً��߆�㲨\܋�E��"��!��3�}`n�*��f�6�<lSh�eJ*�aD+�(ʠ�i���q
1�vy�k�SvܖP�
���R�����,	���mQQ�����v����a�`��)�CT��(��;�"]��]+��[�wێ�Gט��I�mOv	jVAΟ�%����H���+x6�F�k ��fwB�C�ψ�/7ꡲ�����@E�X� G�L;)����L��� ;ߘ�K+��Ϋ����x6�i�����e}��l(
H�-#3��1��;׬^�ۻ��x)[0S�/��>��%�ߒ�=�����1���ٴ��_�c%J��ݎ�����g�U��gieI��79����B�l'R��F
$�>�B��I����ڧ,
��m�����f�)l��Y~�%��4�K�#���/֕�Pl� �}F��q'dl&`�,���m�6�V����5���i��@t���#�.h/�A7#
}6�꓄B.:&���MKX�����c*�L�%��ǟ�dFs�"�1�;5k���[��6E�fy!����뼴v��0��,#�@3c���,��7w����1�GO�2n��*���/�,�+�-����4�7��Y����~�L��r{��lYa$��p�"��g�=oZk�$s��؍�gU��\_���q�K�qD�g9��r�S?��g.�E-O��q�-R�������6�Wdo,jh�9~XY2Ig:1>��3v-�kю��i�yV5���@Y�bJ�/�A/Ǿ���P`&�l����
���]�D(%�W��`��: !�-��/v-��r �;��`���Q�I���ô�W��@�}�#)Zv/89\�����7o�AhOS���Qora�#6֓�vɰz~�����\�v�8���
l�W�?
:��M?�zX����
cS9���q�� �0	
p��Ƽ�icV` �Xk9��{�z��U{�սv�i�.���t(8�h��vG�o}�('kpB��^�B�����]	$�[����p�S(_�Mʱ����D����#�3���(ۿ�*k��kh�j���MiR���Gv`�-*��w����`�u�����f\��T(ȬR2I�ƚ���VΟ-�_y��I����	�d~��^$"���:�����c�0�����8v�4=,��qޚ3�Y��������a��[���J��u�������Gֺ)\�j�ewǷ�*`��)N���S;k������ R+�0�:�>����#�&O!�.@���{pYQ����L��*����|�Z��:A�B���7���I�n�ɉ#�e���!�&�h����Ԗ���{��m�Kz�B"o�ԯ�V�p�U�㸯�7s~IkF�E������DL*�,�8v�Q��?G�d�2���@^hGnȜ�cfU�a(�rR��2�H��[߲���b�
�t��D6����3R��v��Lς��@4؇�3P
��Пꌐ<��l�^ϫ+T���q����K���#5*��}L=��n$v'�ceeZ�\�|vI&E׺��s�ABu�A���*W3��h��[~�PY�q�)M����!MCI74$�����{��ʮV�Hh�\��$�ٳ����5��^����A�w{�-t� o��G�=@���dP[���Z�>ґ��&��T���o�6v�-$��a*�{
1g�L�{A�MB-`%[7��q�|�ݷ��DɝMa:cs?f��/��m������r�Gm���:L�y�p���l��$ƻ��Ƿ��y���! <�7�4��ߧ*�J���0W�	���i�W����%mh?������	�X&��#���z��������/c���3ف��G`��jm��To�44sUm��T|�E�s
�f�b/�0��i,��%�<G`�v&?���-y�dR���#nōA��Նс�^������9��'�����H[��ײ��D&|�x�tO��aDl����ㆅ�[���P
�uN��)���}"�ٜ�
Ȣ�ُw3����c��@�1)nU�W4�ˆ�3�7�dBu�Z�������U�|����������_8g�kٸ�f<.��^��-��BQyB�zOzA�Υ�D�\�k�]��i"��K�qj�OD���c�L�?�s�S�t��(�ǵt�lq`v3� UW��(��r��� ���!/��T
n!z�|���'��r��3�8s������E_���<O�lشg+�v� ��3��P��<lT{�9�jL��v+G��e�U`:=Rw�P�VR�O��-�J"%���]� �	>���y���o9Q��|ΩSb3Pw����2�?��-�d����t������i�ٯ��I�ߢ(s]�(Ri�uڗj��*�C��l��w!�*�߲:˱�~F 'kҜ�6i���>�7��(�Й���B�5��Z^#j(AL�^Xdn���ϱ��y�������-Lp�Q(��J�h�씅˶ڝ�
%m��i�N�[u'���j����_ݿ)�������i��6r.B��sa1*�*
xWO5"ŏ.V�86.>\`W�y��i����q5˽L���3m�^(zW$5���J巕>����s�殻T1It	�'�L:%�BG�x .Z �fID���	>�����c	�s]�y^�B,;#����TR�$�����6��u�����N3����>ԱV��H�)08M�@[͘�-�F�!��P��,���4�!�YϜ#��!i��O�l�ש2��� G6 !����q��@��C-"��(����F@箂�����[f�!R
��1�dq����8f�܌ȥc�55j=6�к�xM꾡�N>����o	̽�b�g��8���}n���x�"`Y߀�'�b�Z�G�V�g��8Й��)������9W�d!Z%���Jy'�j�G�nX�Kzh���㞠�H���5'�I��<�ǚ�u��We�H|#1�R���T�1�����8���6��m�|(�rS�=��gZ��t�����(I7g��uJ;�X)k�l�������,=���R�Shi	ͼ҆9~�F@ۭ��!i�OO|�^��/WC�Mb/d�w1a�k��	�U_�Ӆ[��H��|��MD�2y�x��~tÐ�6�9��b��g�$��R�'�-�D�e5�s�l�Ѓ��h'��&������.(��R	ݘ�[ [����/���4�;�O;v��@��O|�xӀ�ty�,Þ�{hM�Ο�.�v����8zA�m$7ZL��*ْ]���}g�A�2\��[�	ߍ�q%����"����������GR>,ʥ����sv.���]�<8)~��åwEc:���.�V�홠����!��F��/.ݣ^&�yF�c��i�<5m�M�=1>Qu9����Ĳ.{B�%�n����բ��;���˓�4W9D�_=�w�h�o$�>#���T��,��e�{��j�Z2k���QJR2!d�L����J�����~�}荙j�"��؝�A��(E��i�>��->օ��*��P	��1���x���VH��D<�j]�࠵�ѱ0+�ū���rз�)�PVI8��~�X�_�sܱ���X�4���/hhۿ�^��*�����#ZL������	[c���(g��A�.�T��g*c^Q��
7�|�t���{B�/zf~Or�>�$8�
V�ꈰn�N���;�)ݣ��t���~c��=���C(���L5ki�8��2�N�=�����H�c8�oW�t�}z^���z��E>&�H��R8%�� F��	iuqF�VÃ� !��[H�i�vń/w��Y�I�/ØR�����_V�N6��"��	4M�g��r��gdF� �%9L�*�^�浊��Q*�n�8�1�$C�|" @��(6�RH�gQo�Dt9�K��X��}��9N�t�CJq�-�NJ̍0�.�� �噔��A�Ht�`�p��=�v��&�+���WjP}�g
¹t��$�z���	� �m9��y�Ux˨�[�P�te��ϑ�:n�O�D���L��A�I��oK)Ł�ow�g^^�� D��-� H"5v�ӫ��	���k,���%���oD���{������o�Oe�)�+��Z���a�}�����x��FsY.��<q�8�s{Y]��7mZC�De�ſ�l>�,����@��*ԇ�X��v�8�+6Md1��.
��*c�?��R����F1�N�<�����|0U����.�4�C��\f�U;T���y����j��?P�MO�,�q}n���E�0D�x����$����>d�_�gXx�ƧP!g�(�#C�iS"�q:A�.r`�EW* ���X�Q���Jf�q�֎���)��������t��3���N�E�A��ő�����4�����k�.֚mt��xJ9i�!i5��6{�@Av�tb���1u��bʈM���,�9����m��^����[b�m�4��57��|q�?~�Z�
��&?����M�Ј�$��"�2����IT�U1[R��a�KAdayʌ�eré�Γ(+����o��y����n�����	^X�־P�z �%�����O/K3Q�f�ǂl�ZrKJ�[���~̈֒�z*�^y��T>����PZ�!E��@��?ךFJ=�Yer��QȘ.w|Nb��T�(䪬��*�֒U�9�!VD-*%u�hZJ�Dn?��D���x���ZFLf��/do�вZ��+��<�>�S#f��l�-�L�~�e����+������\+�nqn��0eM��`#����Yl�ϣ&X�8�Sc��I���G��hy���g�}�@%���a��2pX��,����6�X����ƾ�����Ӂ������� �󂳥���%��$׆$UqłC��)��A>��zC��̷�@�ePq���DH�'�C�B��������Jw�%��FZ�D�G�<�v��Д�!�6���_^$ �bM�͗����[K���'k�]͜���䤏0��t�+�C���/��P��+鴹C�.�M{���W1����Y-��G7X�Q��(��G�z�(�t��Z�Dlg�g�UEr�6��5�x���V#�P:J��:���亖|b��uL�+Lķ�"�xr�V��o�9�,ّ�ޡd)H�����x!�*q�=�#�ovl����@���)���/���Ɲ'�����V/���F��_럙ˊ�W�4��y���^;P;��gHn^C�C}Ox���[��i���ӿw�PM��Zk�4�O�g���<+�G����Fu�뎂��܌�2lT�7���dJ��T�c��=���S�ɿ��=����f+�}�ul��_�6����_���墥+`�v2Z-?@�z����o�F>y��������2j��B@��ؘݳ�+̧�<'��H�R��N����[>Kh�:��xX4T+欳E�<��B�q�䒛dL�ߒ�GS�(Ez�z��+�π��$�83��g��v���L�9�H68�oT���](k���Ku<:6��	��EIl��fv�%M��Bs/5��nựL�;X�=�����~��H��c�o���-����?�S�{�[�ϕ'��8���P��B�[6��iZ&$����Y_�`��	�ɴ��KkG�.AÀ�]�h�Fߑ�->3��d/o���׽��4��I�!��	���p�o�uaK{� c��q*��f_I�J��e�H����h�w
9T�����œ��q�B�����8FT��zy0ZZ�ÊN�\Q3z*�Y��E��2���*��^ Z!*� ���^�=A�0"76��f�����d��N�;���fc�ZV]��I���oMN���^�=ï(���m3M�/�s����7����������Qze��z)�$�z���U����!A�q�Ek${-�au�a�BXT��G�,u%�t}ѳаބy��SB(rw�h?��O�1T��M�����w|��_���PB������f	C[�{߱=I��[�3���(Dr�7,���W��k���n�N���hv���l�/M�塥�T�(���T�璦���v;f�3��VSD�uJ���s��~���Z��憂{�y�I��Mvh�����On��s��O!���8�зeQ����͍���<yȿ�Hb�� 
0�9 ���&�[���\��`��N�6��;���]�����3I��,l�f��x�ہm
�F����8	�@���7�ﵳ��d�ANU�Sԣ��?��o���-ץ���	q[:���
�в���T<�h�1��3����H����_	)�0h� �v�ӎ��7l%���_i�Ych�$��b��x�?>N�	�TV�f�g�r�;���Lh?�y[����-]+|��z�!@�"�,��WY�s� �E��9e�ꌘ�DB3�r]��h�c^�4�V��F���(j�+V񘖢���j��Fkrq��If���!���ʘ���Nc�A7�^�����/�8�:c��M��}�1#���A�Fz�I[6��bΙ�s�4��+�#�����"�I<�ؗR�]�ԏ\".9�ږ�����������tI|/�~i� ���O�(�rt<>A��P�0֙���{�ύy)�����-'G=���W�4@an`i9��O|5	�]t�U�j\#����ۣ}�OkjqimA���+���vy/A�[3��wm^-�Y=����N�l���ѽU����������g<���ʼ��U)�uc\+m<���y�����B\*��퉕-�x�RyO;�m���mYftu��H�(�W����.ܤ�'YĤ��%�� M	v#}��'P��OFV�*�� �@�rg}9�6_�y9�t�n�	�A��U�Х�Nl����Ӏ�nHvK�.Hx(�1��z��%D���\-w�A:e�<�R���K����G���hj����C���u�LԆ�*�˃��
��3�:r�?d�c���ެ~��s~�������Bg ���w��8t(��*r���R6�<�Yx�I��R�V۬��:��[	�.}�nv�����6���F�o������^�ҥ���>���o��3�O�$��t;,%�| ��ǌؙ�kfj���9b�d�U�7I��c'�AK����t=74�m[3o��B��2(�˜��dE��G^#en��l����q���d`!N I�V��ߝ��:虌�'K��[ä���G����s��a-�C<�(r�ْ�Z'��@��/��1�ϫN���zt��C�\��1�Z�~I�	`�s�	j�9=-�3q��%���wX�s��|�(�fa������7{�y�C�;��C�hs4���ȡᅽcU!�ф�}����6�����p6�j���=?��1dn*t��@�2V�����! ���T�DؾN՝�ƚ�QE�+�2a�-	���^��<�LE��`Q��F�̬Oɴ�	=ٿ�z?r��X�zSk�y��EΦ�:"��mR��4����1�� ?����T$�B���I5 c�	��+�Ϟ$��t# ����V~ud��CË7�hE�xr��v��lo�{1$� ���W�8b�V8�סL���+��r�����C�mZg/���?�Ç�ڬo�K G�}�lb�Ge(�3XϏ���f��7�sJ�ϳ����,B�Z����K�C�^�ys�%fK�6j%��hz�W�Z�!�>Xg��f����q���J� ��6�e�KA��S�cu��ͺ���ց︱w���O�Gǥ�l.�G�qg ?��>`{�&��UFg�ȯJ�6�R��Ǧ��ЧP�g��|n�DI~a�No�r��R݁���.a�s�wm��y�Va���Q��mX�R��W����i��;{A���<�u�uD��g{�vM �TF�r����]�Aj�9jrR|�O��L�q���dPRGm�V��-���#��ج�{&��g�X8�.t�h)�$�-��h�n��*�hDVn�k���yr� �TWCl��-�����/]Z���Pfm�`��e��"k�?*<>��{[��H��o�wyN�|e�6�R����Jw���x�B�1��b����ş�(�݅^D.9��K�Pv�S֠�E�s��.�$���xU��k|��� ��)���.�k!���'��t"�����SÀΌ���������/���4ǂ�D�V,ejZ2�L ���Ƅ�+2�g,*�{�)?-i�rTr��YsgL""��w>�4"�G�u�I�5eo����:U7��vt�˰�BA^����c�MRk��;�X� 1⧮��k��ƥ'��g�n�tylrٝ�~�cT�&y9�_ ����1:q�2�R!vոi:B���_�
��HT`.�õ2�z��v4O�1�N��u�^,Ϲ}c&�&8�\��I�mC�C��m~{B-#MEVD�(�#T7P�0f� �罎���I��E���a�v���7��S�B���5�正���}x����H�H��z6����;��-V���X�6���<C��o������aB��#@Ӊ1�D��O�%B DF�hՇ"��(f�`9��~~bVX�kE��TG�י�S�`�vGo,�+�(9n=���!���z��<�:�Y.�3�+Z3e!����mov�L�J�GB:Y������ܦx��!�xg<��}>���R[Ό�1�c��T\;L�a��1}Ow\W�|3�~"A�x�*�����x&`���_�^�	# dC���`����:`�	��:�߹_�(�*T��r��d���t�Z{X�&r/O"����6���t�ZD�F���!]`[��8����xU���t�K�,W��t��e��.�eM�FT����ޱ���:v"���o[���������N�=��c]��j���\����R��N���������O�ﲘ��BL�YS���c5f�x4�q/)�G�ͨ�c�GU�N�]�F�,Wg���z���؜^��Q�%�`�Hl_���T�f{�W��1R�A$�čj,66ܔj ����#�n���y� �E���y�R	��@��vB�J�E��/�A[j��v�2���~Sn]�ƺ3�ۻ(���q�x
a�KB`�(��#sr�\��RQq]p�m�C�o�B}[h}�[[qQ�����MV��1{7`B��N4�����������\�yrW �~a���u���6`Z���~|��|��En���R�JK;h���"|=�f�2,A���W�"
��Y#�������h38�XX ��m[�7\Ĩ3��V����qT�+�2,��Y�I�C��:	�ݢ�Q��b楓^�JXXK�= $b�uZׅ8���hV>���Ew�Z8uˮ�[�����wL��='s4�`���T�kR#Jj2���;�6���5E�L �^�D��0�$�@Mf�:k���z�W�qM��(���}�NS��7��&���;� x��5f!�@{�a�H�_�ʈ��5&V	@&\�$�*g`�+i�����g����#�q���=V��QE;~e5�W �yHQ�u��W���T�?DN�JkEH�V_F�D�SebqV
��Q�;����5��U������6':��ڊ��jI'S���kR���Q��� 1��Aϴ�l�A��yXzoz��bK")���g%u�|8��q�oWY�dX��z�E��bh�ם[����@�`�{��<p�φ:N��b^9=(Ԅ	'	q~�̢����R@��|���4������>�E]�N�@d
�,n���٦����ަ�F>0�����{xi�,�'EO��ab���m	��$�0�b�͘&��H�C`�d�ړ�:�YL(@Z����:I^��+ w���[���*���[�(ͮ�G��m�/̨�U����Z5 �>��iƲ?�����P�������J����Y,�#�Q����;5�m�w���'>�g�>c�=��J�mѕh��scq�i�J�uQO���z���݉B..�L��-�0;Qn�qɻ��B�Ў�uF81T�# ''򨖊��X�������<�	�y�y��D"):k
#'��s�s�N�V�OE7��4ޅh�poʐ����o���Tz����j���f����"��R����aO��{4�L�$�a�OM*NC���)���.B���/,�@�����
���.S�������@	���K%��������	�3o`1oG����!U�RU�<?���-6$�ڑQiS�̤�|A{�x9��n��/|���0�m�0i��q�ŕ���/	��o㵎����8��t{��j9�tV��<P���,E xa!%�^�L��F�
��;*T��JN���Ӌ��y<��|�V���r5�1��%"�5X�ǂ
�be@1�`�}��v����C���@�~��_krD��:F@H����h�҉MV��-4|%G�r�a�G3a_NR����W,� �Ηa�ba�qS4wa�j�]���M�X�XF.?c����&�bT����p�mCxzk�,�<�������	4��N}�q7�l&���Ρ��8&��G�Q�W��\�!����$�X�qۉtV����(��4ɣ�C�c�3��|3N(t�&�7����4u64�z;ܲ�rs�8v�T�� �2�æf[���r�K�7�h6Tލ����Ò5�Ko��,����7�ɝj�a� Z�	�6�U8�ԯ��)��j�j�]��f���ڽq�K'h�����{x�!�{G���ail������+3�exa��2�awo>W"�B=�����x�5�C;�{~���[��5|�J��y��}ɺ%K�hSM��=1%��7���f���<��Yu�i<�1-�����(#��$+mr���_2��H�g�ų̩OK��>^�.�\��s7e���l���#�Zr�?P]�}�Qѷ3H+��?3��z��7��=�4��uw��9������H�Ej/k�.�����d��,d�b~�1~�ϣ�H�l����Rb��_�/:$��ڐ����߼�KΣ)���S�D�xhe�tJ `'K���� P����5����=�<>�>26�|q�ı�jAd���5$(&����ܬ-�!�K�~��m|�Oi�ʤj�t�ԪL�eS���4dS�g��b ]��т9��.g�
�zC�X�+��e�$Z�I�.B`�k��%-�`�Y(�̳�$�{X�����G�`h�.� �A
�a~��(%jÿ5X�7���r� �rS��J9��hS���B'%q��!�(l�xrj��Q��-�:P4.jѸ�׮fv5����	Ħ�5km��mr��ċ���Q0d�y0�"�<d��"�6w�h�d�����^m���>��ˣ����0��v�U�t��(}�1�q���m`�nP�3�!�p���uV�v|�3v����lS�|�jv�O�K�� HYY$l4�u�'6
~��,�X�;mk�-:�	��IB"o5Os��T��)`�� �n4s��t�.��>�se����)���ۏγ?.��,�
���$��A5��*��C���qߩ�H_�O�$=�:��6��"R�G��t�u8��bS�fl,Z�09��Cў���߸��	4����|>�k���Ɔ
�u�ŧ��vu��Fէ�"h��F,dڗzPs	{;�$5U��JT[�@��b������v�3Ӥ��t�G^�!��F{Le�o'?qN܃a[��8�z��74;e_�w����.��`�5���AI\�+��똯s���q�..��g��mJÍ���;�; ��f_��o ,p�$�Ͼ�֗���e���K��Nms����D��XW�O��d��E��2|��.�����?!����x��3�0�vʬZ����F�b��������b0�*G	)��KR��"O�hwf�1խiU���Y2ᤎ�>}����\C����>�E�VD&��<?Z[�l�Sc�v��\�!�@9��Vn�_��U��>T��n�*��<ߜ�Xe�g��_,�4Aܜ�%�(���f���4r=�'FNN��ɫ���[ g�#p�֔Y�A/���B�c����s��A���(gMZ�L/��� �j;��
x���n���n ˠ�Y-0��7R��ۥ=A5�;Wx��T�g}��]�Ϭ�{��h����N7�j�[�,�^���MK�=	����;�!o�W�߁���pW0�2/��e����N؇u��6��_y#%��e��	�	4�$dx&��%�h7��#X���f�
�oXD�t3���`gb���x�,	���;v�>��P���j�I��
Y�g��24���m%Mj�w�����5��/QлMw���Z���!�&KĐgO���:���BB�ldB���*zWcD��u�k��V�tUn�Y�/��<R�P��'�UєQ��t�N��4*���􈹑�Y�͊�jsG�:Np�e�a�h��9��3O
�S�r������ts�SB}w%L�����lsЃ�Ka�ľ*��l=���Q�
���V[�<��|fj��І�u*Üc�7}J3ȫ�JS�U2nҐ5�����rk͋\��wx��y�M��c�zt����D�������Tv�{�f��d���Bʳu�[�����.I��qkB����-�5R2���h��m�	�Y�69�dd�K�~�r3q!#�����5Į`�,�[��YD��A���Fi���	���<�^�C�F���J+yo��B�|f��'(pr8�-y�S$YM-���vbHΗ���p��	��`Vn��� 6�0jy�8����:��|O�D�m�3��5}�_r��D���2_>g�[�
�2_�Es��N,ަ�ɊR�w*�4�ݏ�v_��5��2(X8��tkͅ�dH7cb��Tµ1:�x]�f��t�h*�$�O��S/�c��:�jh�����F�&�/��l�����=	�re��5�t�!K�FK�.\h�q'���(Xja�z�w�+�D�p\T]��rjoEVXe
��	֑)R@����V%,�dJl����1��N�
^fG׿������7e�
On�����]��B�4CV(�N�p/��EqJ��U;"�䩜:�������sD�ycl1�X�LH�[��hOdͳ8ȊQ�����s|X<��4��,U����{�ϋ)�g�A�|3� E]:�z3��td��A��u#�o{@"甛�)����o������+;
�f���]��7������yX�,�d�P3�qXws�=W���M1$c�����j-$A'��a{��@�Njo!f���>����q��]o����#�T�I���+��b�pJ�5����Z���y�͚��T!�_	�灊�R1cT�'2擨�H.�툭#CA�[�%����k��2�j�Z<�P%��O`�\/=��5{f����:a!��U�����D��x��v�[�� ����DfK'��9��%��60`��$a�b�"����Q�����6��W3`5E��~6�2�QkB�g�q	+���
�;<��-Y��=�nY���ʭ�q$a��&t�tE�^-\�����$��
�l�z6��!\f8Ž�3~99̌�_�|�n�G?yK
`�a��h��6n�k�ej�I �;jb�HcQ"*��-�����"�m�f��}=�^ӗ�b�k�Y�W$j��\��+?���)�����G󄇛�{�s���^�B�=�c�$J���L��UH�B���`�Y+{&�eR�Z��wN_Y=r���6Sq_?�A�3O72���2X��-��5�u�*����M��lc�rv�H��LP8���S��3�m���+�y�q�Pl�qo�F�t�_H*i�{�.��V�KF<h�9sJ��F"�-|-���[W�a�<�60�����kz�ᅟ��L���r%�샽��J\���d�E��I9��+Gw�ؗb��TF*��;��-�l��ŷN��n�q:�݃ZѣAE�s�	hIU��"M�0�J��C��2~�k�P�����F�3 �U�3���c�}����n-�?�*XC#�dExZi��NK,"�����="�����̟m�M9�4'�(��G%订��U�ƅ ������S����f5�EG��%h~Oy�u=c��w���P��U�^M���ȭCU�@�aa��� ��}IDV��b��$�3ǯJ��� ����sU�c��?Y|u!�Z�;ld�} �]�rdҬ���&`�5���0���cBF�R�����P3)W�O�<S]WB����T���(]����.���B�u���1Y3��zQre �*�Y�����(S�t>t� �[�͘�tjI¥/�D/���{���H�=�T����U�.�ZKך���Yp|��g<����o���Y-%���lvD��`jjD���$Wu��T����32sO��NZF��YG[�.թ)��:��iP5 6��b��\?���~ױ)Z�ړ�)9.8Y<��a���7ȧ-�9�H���@gg�v�Ԃ�H s(<�"��op%u�4�'p#_��*���<��M���>�2���)���)>
�z0�"� ��=�����O� �T�Bv" uk�\Uz�aІ�IGf�6�z�e����6�8j�c��1#���}է0q���B��I�n�.�g�<�c�֌�tjz�n�(�>n��Ԁ,
F�3��-l��#Ǔ�M񺀶k���
h���Z�g��������T��^l����\��JM���V��a�� }�G�Ԑ0��s��`�m�����_�t!V@�)�M
%�L���*��;/rTN(m���9 s}4,N�>��,�Of�$3Z�
,�\��d̼�,�Y�aS<�Ǻ	�$Ց��97r�	�v�!���r0?�b�ߐ�}L*6���35��M�8������+5���%���������,[���h����3^��!\��MN4�\8'�z��f]�d*�n(TV
�c�6@�Lĳ����J#@+���K�Dl���^�)���Ǯ'���O�v���M�Hp"���gu�Bu��>s�?Mc0��$��G/4P�dJ&��l�\�7,��0B˿0~D�:�i�������q�U��k�F䰠n����(/z�5�D?:g�TMohy�9� 2�'�M�_���q�֏�w���΄�;3�[}\�������[�@�b;Q�����.il�@������ځ���N9�O!��-�|��)�v~�8O���G�x2��o��#8��d�{�1Љ��Ӈ�}0�wd�!qN��|�kϖTH�|HMB���.|�� �_�3U�bւN��3�Ǔ�!CC��n�,HM.��9@�|�N$����y��v��/c�-�Q�˛�d������^�aQ��W��@�1*V�s�Q%��f����2���m�@B-ޖ�}�b�|}[�͢�,�N':9��0$�����*��u�J�yl|c����>	��9�3��K7m��g�R�	��U�!�Px ?���)�T��&+�2X�����jf��^*�}ؓi�ܙ��A� F�q*H���B�-�����CP_�2�́��DjyG���L���S�H�i	�{�~�1�\`�)-�����U� �Y	]1M��ZJT���r�Ń>'�(䊍��D.�$u�����WX�4���D��K�s��1�Y��ꨖp\\��U��`Q�z�@x�/�+�yG'��.6����#�YWKML貭�0���<ma஻�P@>v�?��YIF7�c�>.]Ɂ}�i��֣��Db�GP0�|�o�%:�6(�!�BX��� `6�^�ǚ2��rHY��b��Ջ�T1l���>�ȩ� ⌭8����A�,���;J0���W|�^"e/BQf=H�nQ��d^'�9�����@&-<�]�o����G��٦8��
��,2�9�q�� ЭƄa����
S����p^#p�y�
�=���q^�t?eO��X:}�ҥ_|��dvL����9�e[g⏶�}y�kWaKd0֘KğO�"�6�PkC��J�#R���I-��;�.��9����qd�wc,(�Ϳ}��' �����Hp��=��F1�*(M7`�F~�g^����=��8�b�1;����	���m9�� \����x�9�R֝}��emf���7�
8���O�ߔ~2X���X�|Yd���
 ���A� 4˫�����H!ͨYC3枇�>��q����!�<�o���D���S�jɱK\J��w�E�N��԰Ȉ��M����+~�x��1jiTl�RE�.����n���'���QE�I˵mT@[�Z0bL���o塌S�{�p����������k��c�a�M�qP<��-��Vq�R�9ӷ=�-��'�2��1g���j����&e�&���|ZӐ��O<���T90�&l|�`��������Ņ	�+�.� Ϻ|Ն�CRx���-���X�:�l2�Ο�Y&Ϧ]R��H� ��E�e�,��x�'�k��p>��<§F��i�'��ֽ�*T���B+�_g�_ô��S����3������+x�o��OF0kLߐEo�;����(����4�\{¢� ��R,�����3\+�<�(I�R�)P
���	a`�8�k$D�m�z�z�%+�I'?:����D�'�m��5��`)�~���Rz����}��{T���X<�����#]���-n�$�s��,;���z�~��� �ұ�h�(�^�$(�uE��/2E�d28�VW�v����ܒ��J���d����IG��4�S?���	/E?�r1|��Ig���Md_�T�Vb��Ֆ,���w�ݹ^9nIT>!�I��\��~�����E"{m��>+����܅>(� w�+���
�x��q��h�J���T��?]0���j̨e���NOz]����o��MQ�{������Ŀ4H��؀E������Pu�\X�����������
�����_A!���%쥵�On
=G��o���_Epp�P���g����a8&���\����y�k���Yh�X���������[5�!l��YS�.#Y�V��rN�A2P�ۀiDv];`��.����_��>�/�[%�[v\�U�H�+��pa�J��9+�*5��J#)R���7`-pi�t���	��wc��o����PP�D�u��ݖ�`���pSsǱ?����Q��~cD`,�ʽn=e�)H-��L�̓;�V��ob�= �����M��۳S�JV.ηL��8�t�e���=��g��wݍw"<�G�O�U��.�CC���CY��fb��`Bf�����z$*{�[#�1��1��ݽ�E�u0���P�k�����Kh�0J1A�I���'�r�8��Џ0V�*'�F�8�-,14>+[����d}Ø5^�FH��3���?&����ة�9;M_��- �>����D�vjYJ���a����֝�P�P�a(3s�\ﴩf���sΧ������1����!� �������y�ӵ�3�M2�R�گlE�>�-���_��I��݅bLA�`��F�	�m��V��'��Y�����"-�k.Nط�Ů_˯1�-x�%�[t����8��k�䬯���
o����b����u�QW=�;����y[�&�)��%�Brc��ӬH�_y#Б���z�-M�s#��&@[����k���.F�s3�6��gg�!���pc�	ͬ��!�b���+��M�p4��A^�VK�ܪ'��F����EѝIP�b4����_��a�U��Ę��Z*sx��EF&ˁ�1�����x7�qΉP�fS��b�7�#�+��<q���n!���/V�Ǹͷ�B�/��cjk�qi�*��q;T.��/W��so���'�!k���7�An��������:�yPx����e�4���J����w�@��\R��6��b[O ��&1�h6�U�H���{�KN �� f�Ł�L�
)	����wP{��&''��b��mYR��=��F�a1��9_�	�%r=E�2E�[���(����t��$���h��V�(�0���d��u/����{��@+�l�a�)���U��8�G������Y��@��IM�u�KjQ
b��0�|����]�=4%+BR뗭��%|����	�NC�m����r�e��!�6�p��~q#���`�����g�6+H~~z�P�0��\8?���չ�tKG�_�\ӧ�hr���7���;�'H���&�8N�~��a�����x���T�����i[���d�.�ҟ[�<9R��A�B�/>5�nS��UF��h\��F��q?�ߩa:z#�=��k$ϊ�u���5/�B���ˤ����"�?X�t�bY@*����7���a'����*ij%��+�R ��o��1��H�І�խ-6�W�?!��6���I�&c��+ˑ̭����]Ԣt���R���������u���@IR��i���qE�s�m�E5�F:r�A+ ��3
:����~���)ř�P@S�y���.�i3w�6��}XM��Ĺ����*��[��5�n�x���E�T�����ʹ�Ӻ��l��/S��}^�7�8I�)���sY-~c!�p��+�ad��U�Ä�T��b�ܹ(ijЍl(,�K"G���A[7YC-b��1Q$�׀��b�[8�)����d��ш�)��b*:b~���5!6��g�O%-u}gڡt ,ň�E\�K��c oWK���&��u�n�Nz��J�|�G�u��b�궷���ݿ�(���g������]��O ��u
\y3�G9q�Zn���t��d�Qq#��(�$V�傀^�P�c��&��A��>�ɺ<Q�	�Z��O?&��1>x	����+!ڥ�;��r~D#$��9ڔ��F��z��B,�G l4��x)��K�7��-]�/��*w'z�O=��u	��P���P�p¯+��)���6���tY�# iZ�]���]`"i�43�3ڳ����hɫjC`���K��({8�c#=[�P����Y*�������3I�yy�Q�%���
(yyӎ\H���)��u,1�C�b1�JzLr)4D��=w�
hC�T�Z�q� *�E�U�NӼ�{�[�3_X0��/���>bT���#	�yR���I[uR��T@)~"�3�X�Љ=�c���@UL!,|��%�� ��Ks�-���8�`x�DA���U]����Q ��?�>���|`CsLk�[��=���O����D̩[a��c;Pl�o;$��R3�*h ��G����ފ}�/,2 Ҏ��dk��p	݃�=�і�4��f�a��A�6	���%���j��n���QJ��ֽ46<��+d�M���]6��:���&�!�D-".e�ɹ��R�V<�l���-ܵ����sM~��^\F�+;\.U������ź�h9�ZN�Gnڛ�kp�>��(j�h�P�d�i8�>ݘfר��G8�^R�!��Z�_����?w(�uZS�R�<+\J�\Wq��l�Yט�I=:tY�������boo�Y�wf�i�nT�`��8�v��M��D�&^���"˺�j&\ ��ؑKJz��� 

0y��.L%��8f:�����
(�-}�dK.X�L�Lj�����Н�����q��1���?��Z��������L㍽�e}W������X�L���ϩ��I]�HJ+wz��ҏK�z�W՗Z�}�X"ϰ+���%�+h:d%�3�ړ�?�
�ۈ&!!/f��uZF%g������
�'S<����N��EH2��T�ߞ�ܔ�G���7�o\6^������S	�߃�}�K��Bv�Rlm�~��Ņw�F��f�E{P$`��e�J���j|�Q�/�ˆl/��~8�xs��	QM����\�""zV�g)�r�Uc&�Ym9�QdO6�a*��@3ʟ��˖Y�$��	ut�õ�=��S�����I�~�Ig/q���p���?wͰ3�}�ѳ�TP�u��3�V��E���)N��⺾z^�.���X���q�����8����ǥ������i+���2��^��C�(���y_���X6�~��!��2x%snh�H�|�H�:�ص8�.�&�rx
"h�"��z��Agj!o�"�8 ���V�� ��	%F���Z#lȞ^���@\�ʇ��kɢ]�Z��w�j�U[K��H�Z�l5�;���= (
�,�Vˠ���]��ՙ��l�lQ"=f��=7ݝ�K���Q7p����dC�5-�xR�i'-6F'��9H��S�(̞w�e�(�5��֦|ֵ�F��z�(\\�V�Km�������U���蟋�?Џ�u����&��CK�h��-��ئ��͌r�3�e�4�K^�4�J�5]W»����_���N��Kg��]�wuEt����)��Kv�Y�F'\�+��4�z�U|�&�Rv�s
�"и��A�����sX�����1���.4vz5�Ә������q]|@<�(�9��A�k���\�n�X�bq�D+�r�9��Ǿ��#WUY5ӶB��O%ua�W��yi�2���I�#ݠI�ܬ��T��&[�4/����t��b�䈱���vsdLtq��B�g�F��T� �1� �?ژ��9�.���oe��,��\�+��CY%T���Н�%�B�!DWլ�8~�q�op<����i4���ۯ�V���	���(���$UY�X0E�췛_��2ן�\�>�F�V��y4�f�s:��"�rq�׎��ͯYg���{qo@���{�e���%hpK- A��"q8,Q4�wMٝs�U���ᝪ/CS�U9ZR����D���_c���=����	�1K�s���'[<��ؽ#^�ܸ�ފȩHj�N挾͗������70ۿ��Xp�ݜ�R<�h�I+��G���T�6 gӪ�0����:�n�s�5��6~����$�W�(H���j_�R�_8\\s�I�s�X9	�**@� ��!����@�)���B�=R��d?�k3+
Ǡ���XL搓�=�;Y.�'ј��}:u��M�����}ڥ0ٮ���ڬ��������Ql�����8��	>���.�z$�7h]z [O�,�)y/)�u��&r^ɗz�E���f VRոF"p2� �Ӟ�����H毕��*�ҩ ��U��8L7�[��2�����>}	�U�}��D��i���ٸ��j��Q����'!}x^:
�?p&$]����Y��㒘����}�X�YK�=3%��Ĥ`֜f:��������]��G̠]��5H`Xl��˟����F��6�zs���Zb�Ԏ<r���o�Ǫ��KMD��"K�9B��
g"�=�����D������c�=&e��q�m���TW�:�8s/�L�{��%[���`�$}�@Q,�`?�{��J��+�G$y n�����1�E+n ��$��(\�蟭U1�\�D��v�R��x75�do�5��;ۗ�!��h��6�{4���-=ʗ8�'p��g�4N�,������&�J��~3eav��ͣ�}��\��_t�9�g���N(�3�B�B�Bf�ߛ|��f���J��Yd��:��b�(�ұ
��O��X��V>@��+��r>)��[�&�*�hwԭ�[.LO:�#x�`�&2��}P&�d%=7U��%¯c~`�Y|�^��q\j������%��R�^���;�w��0�<�Q:�H�p�\�PPG��U����h.X���H֤؈M"�:�������k�@j�sq>V9/$��K�A�f�)����԰vԹ��3�a���� d�&ۊt$� �S<Tn� ���]Hؓ��4,A��[�e<�0?u}���(ei����q��p#��U��ЙhS�4�R���	2��68�t�~�3E��w ����}b�'���;]��X��%Ȏ�N���y�S����	��Yfd���~l&��Ք��F��0�6d�w�����$����{��e�r�>Y|h�r!!���)U�<�i있����3q��8�Ƭ�R���_��M�a�B�7y<XJ��-Y�4D�1��ؿ��A�"
��h��C�$V��7y��n�t���O��1���C<)yci��z	;V%й9��{��wX�Z�l�9b����A@����Nh�$4���^�vZM���Z2��+3��t'?����8�3Ij�X֖�\B��<�K��/���G�b��9&���DX�I�k�N5'oW �����].}��4aA܃`�Ǆ1�L�=Ü�I[1���
��`]^�|ҺE��ӛ<��:������'�������$�w��y:dd"U��#�|�:��Z�ZC8el�m��Y��!9����� ��/3�� �4�ZZGp��bx;�T��8�X X� �d����X3)��U-3��`k	���A����ۭA�M� +oiV��x�*��ꄁe��"gr���m'F��O�)xd8ܕ1�P�s��=47�P�A���.��Zg��Wޅk1�cFo) ��O�;��&�z�^��x��% �F��̧ ��"���SZ�"uA��w%���m�Jj���I%�oY׌��"ů�*��q��&��9��M�R��k���Q-�9#=W�X8r���$�sM@|U5�8��u-q˿B�����F^MP�ܥ˖�M����N<9)�G���o�~^d�+���0�ʦ�F�Z�L77��g{�T��<[�	?�o���l����3d#K���^xxD����ٰ3l2��&ׁ��p��z$����7;*���@fD>)�����'Z��_B��u@n�P{S 8j۱^f��C�s���v�b�4Oɺ���	�/�h��R�<}r����e�b3���r�8���a�ܷC(x��%
}g�uH�O�4�B�fGx���f��IáK�^����+��6\iy|�i+f���B��2�9�~�7[o5(�w.��(p�eH��v!"��7�5W>?������d�,I@��+'�AI�04��:=�����@����ȥ?���8]O�pts�����zϡD�\���`���r8����1Zbw��W�y����}zrT!:�������;c��x�&���s�9��f'��"�l��ȉ"��h�g���P��"���6eGJ���r�%�<?@�HqSk�U�RǇ+�3w��u��(��O`��X+�Rl�X�)����-�p!_���Y��T�i��C��Ե���t�|-��r�d��v�f3�a�&�kz,��3e\�s+����gDq�ch�5T�x�a��+T���y(��媿"��S�0v�a��a�T�0�������M`�����cb^v�E�� �bg\���6���q��^*~���Y5��0��d�-�XGKGZ���Sv�ы�}24���Y�q76KG�-��ߥ?tT���|dZ4��ѩ�)��D�!�yZ�f��6>kI�F=�:w�A0`� #���yL[��^r?���䚤U2�*�[�wp��b�[����":V�k�ղ�y��T/�܀��<_�#Ņ�ڌ =�ڋ��hf��T ���6{���
=#&`�)$Ra�?d��J!Kc�]�UU��k۸�Z�Y	%]|�FJT�������n�Y��Lsȟ'=�N��+'˗�*ɇ)#3���'�pIu��)O`QU�g���PB�"jإ��*5�c��ݕ4^�L�4)���y��R��&�`%���&�'�薲A(4��sF �0+ww<�i)��%�;�̒l���{���5xE"�ۊ��vi�}9I�kǀ�̘oo*��(W���Ȗ�V��
�����w����d�iI��c������Y���L4I�K�������r9,{�c���[��8`���w��M��O5L�;�(v��Y:�� -e��������K�(���t�X��htZn�iZq�E��Rq���^��|�UJ�F��nf�n�{�+Wc3�G�j)�u���n�I����>G�l�\Gj�Hpd��x����D!��/�좓��-&svG�����B|x�'���ABp�6dΠWrr��A~$`�N��#@��}{����o�)|#�=n"�MSj4%q���`]�KwV��=��T�;��������MN�Q7#A&x�6��ʎa�DN��.	*B�� *`���u��ߴl���
Pf`�Sx���-��/"��X�n��d[a.L��N�R� ]����KI��j���wU ,�Te�,��e��QD���Fu�$�G�N���:p�.�D�ۢ����㞟
���D���8x*����537)7NS!(޻
I��5H�Q��,�i2���}�ٔ�8 3p��3���2�}I�����=�-uO��) 1m?��*f7 ���������^=��H�P]�b��S�����i�>�t�_��IZ�e���˞���`�ϭ��z�H�E���x��J}z�H#k|�b�+=xo�-&DC�A���H"M�hy��ֵ,��"��[�Q�f����3(��_�	�2�f�|o�m�|
�yW����Uj�����V*|�Õ�o6�{�.^�[��_"(������~`ٿ*F���ߝ%��c)Yԋ��YgL0i�ٰ��;(b��c���+�H��}҂�ۄ�J�'��}c���	����[� ��'|���r�-� �(��G�6�ϞW�a��#�K=ד�S�^��T��<�o~���w~@n�"��ז�ֆA";����b{�\^� h>)����-�W�����k<����A��u���7�v���۶��S+���ݻ����L�FG�N��ڰR�x�)���0�]���z�諷CP�T��v�z}C!��R��	_.��'���<f�s��l7��J˽dۡ̅>x%Nt|�h�Vt���U������f����������E*�]9hU�}3�U��w�[?A�+�ɝ���FE�=�o��O�=�G��^�>!aEO�^b�'���erґ;��ݿ/��&�*E�u8c���H�t�l�ɾ��U�Jt��z���׸�������R�Q��Icyr`N��0�h��	��Ia0�r-Jů(���#�őc❡���!��A
�J�N΢�sƞ�.ɉU.Jw]ƹMR�J`�T]��<�g��ڢ��٧����nm�۝������K@�^I2`�C�\��Z�D焐��Fs-\NҡD�y��_s�iMW�Jz�F���!�^ﲜR��̰�#����G��F�����&�7���\=(�����-���u�<�'�Œ2BJ,(�5٘SL��l*��1&� hL�G�!�v�_�A;<����,[̈́^�#�U�1�S�O$L[e��|9ʁR�F��B�̭� 'Ut�O�V�GO����FMQ*���ňh��h��8d����\�IHLG�*�, �/|���~��DC,�e�^!��0M�- `%��(�����P�Iq��v�蘍F4��b?�:X�=�0����I����aO\����A�p���\~~��[G�f���Qї����yi9�Z�f��N5F�-(�<�i	s������X1��^'r��l�����T�q�tGp HbK������̋{oWw;�a�`x
�Q���(iB�|�ar�5�nT8���G|4ҞN �b�,#`�t�-Z��r
��>�
��
�w|�f,"��X\S@Ϡ���>�L�����)i��_i�d���|t����U�d[QփZ�x�9yB��[;�=?d1�C#�+Z��8�����n�Nce�G��ΦR���:� ��I�v��!�Hd�Ob`ia[���Y5a��Q*n}�0�.��4�0���ɭV����hj��cn�l�=��5�v��փq���L}��.J
*��G�H��[u�!o��"��(t��:�Li��dN�J8P�E�)[��`�jV�-2�¤F�`F��}�i��s�U��}�+�g���F-75L70�-��3T������VaT)Xy��7BQA'�x���YiQ4���``�q�H�M�fei�c��s]��[T�E����-��{�rv-�����W 7 ��{; �%�enH�T����Ի�ԫnl	ζ�RÁ�x�����\���g��?M�g ����6��&v����E1����@�B��g��RG��[	�=��u�Ni�U�YT+���p-��*�o%���+����w;�7nO͜�?�+�W=�2�X����{�H|�r�/�UAm23��i�O��G����-� x��9�#t�C�\����Kī@Q��I�{�j�5�����vgʹu\�ų���<�3(��@�D�����Dq�_h�r����K}��Y7!��B�dSD�?P�D琸j�1(�3���[Z��[g>�la92r���#)Ӵ�q����ÄPͥ�e�Ax|���)蜜��iB��8��V��Qb�\���Km�@s�e�p������7�`�,���8��n� x[o�M��q��[ �oi�c�"L�-i�]@d����҆!)�0��Fnu���r���+�Q�nk�w �":�*����S����[��S~d��K+/�h�?���U�^@.��=�b����s�Vb�ɐ�S����υZb����h� �g����6�f-T����1�?�~��5I/��g��C���-4�i@}e�ɛ���(065�_�7h��]2�ml��U��c[�[⦬�*��t���ԍ���Vjt�(�\s�Lɩ�U��o0��?�-�����>�ao]�R�e���*ﺇ�
�8�5d���y3�Tj��T�hBB"�'�	1�d$c�<K��nV�:h3�=��m��#lB��ێnx�0K��X��׊�mp�f��U�Yޯt+�ճ��4%�"7�NeP���ID����_�,~��(��ևa����})(9���y��v<�9E17�G<<��
�h���U�}�j'9�E1u?2��s�W�/'5�u��F����xX�
T�"�%3³���R��ipeaq7�w��h�t谰��Q�9��w��f2��Lf}���ID%�l�G�K)�؈��.�<;�I��

!`"� �4�og�!��6m�$R�ɥ����������	�@��(m�/>�{�#XK�g�/��lt��B��s[��͏����p� x�J��Z���pA:��pKjr�6�� VI��k�d�s�z+e�ϛ��K�D�+Lш'�t�?f���m��8!���l7�e����ǅ�����ZJ�#J���v��`פ�7
�DV*#�U�.����5�.�R��)�ө��?]"��t_�D�%]�0���cFg��:,���"U5n(��Cet47��{��/��=��f�C�"R�1{Ɉ֟Y#q�H�	.��tv���G��A 6��7��e��hi�A���o^�}����T� �S$�}p$��!��ka���.�~��žHn6��B�V���C�)���NrO�4� :\�ݸ�J��ΠFPg.o��`���Dґ��Q�J�rS���b@�W�m?�1P�D|���S|(W�/BP1;��d�6�P�-�q�
$�* !7߂��c��6�kV�Z���w�97�> y3�Lȧ:���mˈ��C[�~��L�&�������n9��)���vM�Jߩ�� (xE@#1�_e��}%/�|��;���kc��d��cܞ�}���c����Cﷸ�4/A��o,���y����ʄکZ5���]"��=�˷�ni�W=�9��EW�#�T��e1ݺU��� E�QU�I�Y�z��Egf<ʜxUX�V��t1F(����3�#�SY��Z�쮀�떇r4���sB�L�}T�8n�$O�J���K%����'5���ѱ�O<D�Pj�K�
��6Zf˭hy�Y��͎-�}]��!�IP+!q�������<pq��м���v[?p�X6����cnx HE����E-/��9�����f��T:HzVr2�w�T�d�S�]a��XVܠ95��ܸ"�z��8����F�[�a���؏J0A���R�C(�m#:"������M��m�3�,A7���46Ί�ŧ�c��AZ�ChS�+��I}�N�<�V�0AAr�8j`H-�o��F-e�md��+�����8�@�m��$����T*�i�-9',ݬï�����a ������3�@5�Z*�s��$y���6��/[2���ڻ��V�^�:V�����x�y��_:e�#g��7��S�y	gVY��I�F^�^�mB�ח��9x� �	!��?�CI}㕑5M���x/�r0�@jMI.����j�R���5Y�ߡ���Oj��l�4K���R(Ӧa��ѕ�3V9�yEU�������u
V�_�L*��$�Xh�M��*�βb���z��x��ײ��K���u�
�������w}����]3�`n$'���+'�4�&��2�~�����$�d���e!<P�m����zd7���_8(qO�����g>N)������DD>��d�N��9��fcj�Rc����������X�o��ٝ�h'���������!�"���iy�ɻ�P����O�s�>��Z����SD8ܧ�����*;�F�:��J��ᒵ����J�<���s����g�.d�>/] q����t=����=!����R<���8Ҧj��S�32�&dE�#���-�t9�*O���5�!9�S#3fY����V��uM��R#�6w:���!��`}v����x�U����w����;�*��(Z�9�G���3���0u�-m!�wm��t� ������
)����Z�|�^�XC�F��H�1����T�(��,h�1Qnk���	�\���DS3�傺^-�40`�h�f�-���&�#���1ԯªt_R#1���0w`����I.��<C$����)�y���nf��ACm�Iw�Y�T"Z�S�U�6jM\����ؤb.�$�Z01�#�~)_��%YxյB�R��\�w�1"����:P����,��V:����{g��5*2�̉����}�E��2y��h��sO�������1Cs�εЀ��")h���5�T�^���o5R��UM�-pk$�z��v"o
f��b��]RB��l+��AuɑGp#�Q�C`��|7�����c1D�-n��\e%cx]��g��2D��XK٠��=��ժ᳐䙧<���G7ccn���aq��"�{��	^����q�Sx\
R5}�4ams�9��/��?��3������m�u[t'�L�#��D�n�;�0��	�BQ"(�)�.����-��  �S����G��]�l6?&Y�k��[�j@����KI���3�t�zs�Ϭiu�d ��3~������C�~�l\v#���U��;5P���]��y���V�ٲ01�G��*3^�@��?c��UT�.E��mj$ȵsqH�-�K��n�+�]󷉛�I�̈́����=1��ë6w�{�v�S�?�*/����w�T�H�(�m�&*h��Hh�͛��O��)ځ�E�|���u��P=����^b^�u����n��kM;1���\Y�|�_�̍ �����
G$����P�Vl=)ȏ�%���W��?f<N�dߖɜ��sxDly�WN����}[Q����O�E���w�-��Z�Px�r�����s��'�Ս����D�B�w�񲒂:���䀏�>�X���}.��W�?ܜ]��C'�r^y-�q��`ܹчv�e֛{AR\���J�kp��sB	SזE�h��*�$�Z	7���nD�2R�-vZ�Q|V/3Λ�U�BH�/M���g��TX�Cq��p����~D{��� ���ܟ�o�
"^x�D��*#)�
�:y%C��w��]�w�h�n���.���
I�!��<ז=X�T�1<�֨v(�*A]
jT|j�KY�v���5���<��J(=����UI��uo%Z�[5c�Ӕk�:��wL(�]�&dBŊ��B�x=��!y���<���^#"���Eku���=���B�Z*�#B�N�fZN,�|�n�k����#�cD֏n �Z��W�9�Xc$C�����w��FgnFN~{|B#�m�q�s?�"�;/�2�@"�k��7�~�0n��8����4w�)��ɕ�|�h ���KL��A-,У�,�Eu�G�=���Ee�z�7���=l&N/����m$����鶌F\Q��ytGcڔ�-�S���0B��]`��p%f��G���af-���S1�Ţ��`E���XTY���Ke$aFm�X�1.��	9��-M�c\�xl.�ß�a#S���1*��Y��`�� 0l[d�����\�ǖ�9?3U��w5�]EPI����B(�{����"��@}��ojc�2c� 	"�Q�a�ᗩ}�A��΀hl�1H�M��Q���x���O�Oj�F�����8�x��h��>�	w��z�z�By�TGZr�s�A�,��Gff����1�����#�piK[� �K��V���q�����%,\�)l���s�+��\��㼤�ӈ�>�t�HT���^۷=nk�E�^&R4]*G�<v`�>�7��ٷ5,Չng�+T��(�w:H���-FP��кM���凬_u���Z����u9-�al��^��L��N`0���O~JGi���v��		�'嫢��ݜ �@��H*���BkMN���*����nH��)���e�~@ńц��>;���|y��0��t�&��@�mZ�C ��o���2H޵��D!{S��9�sJ�+�8u���+���%�UT��ܳB����� �!_|���(^#.���`����;���k�;���W�KIH�#w-)ʆ?��^��,k����Ry�"�k#f�G���EU�����@��!∷�V�[
%d�����#�<h�6iA���Lr�<��uT�uQKë#��n� �`�Tw ]��;��)�V<���&33|I�b.�H&2^�QS�0KHCvp�ez�J�P�d2G�'E��y��O���9�]URD���q�kT�:�\�G��3���R)繯��;\$�Z�O�-�x��%�(L��݂��::U2c�٤��߄u�B��;��#�<��`J��H
WNY��o$��]X*H�	}x����^��1ӓ�8ǔ���q ���#XaO��`#7����6X��ýOզ\�TL~�U�F��a3����7~��S�e��e��#���(e�i`��~��A���ʮ�=�R�K��o\V����fP&g��u�_P�cH�vRI�+bf}ˠIRi^����z����&Xr|w~�)�ޚ=)�f�1�]o�H��`��Di�	c�3j�X0���&�K�1�up@(������B4�q�3G4p����[O�w���`�Ez_M_�o��$-��$��b)rl�f4�����/�v�ϝh�/�@����6j�� `#�G}��Y�J�#sL[�����[�XB�
�A�<}-Y�m�_r��\B�l�����%{^t�R���C�;A����;����SAUzd^�rj�P������g�n�8�}�7����)�����!���a�7����a6e[@���g��~��X��=��3��h>sy]R�#j��F$nJ�dX^o�K�"���2�TT�̣�6�*I��`}Ek$�60_p�i��]�1������3�(w��ј��V�ML�m#_ϲ��ZC��`�V�$�Hީ ��z"��Km�7*kstm/�;���](�T&�[�4Z�tغ>2�H��@u���oR�/��}�ku����0��-���W�h���H�)�ʭ�W7�_O �`ފ+��0���ӧ͓��N��n�O��"}���=��%������tq�Y]��: )wXA��2�X��0�b�ͻ�^v�^��K�٘G��e�r��z��l,�)<��9���#'4�~x~�2 �,����1v�Av�݁'�颈�Ni6Ar+[l%��pn::�k|�����#{z^����6 -��^�Kh.�fo�!Q�䊛B���Rc�PAl��2wa ���_���ٞ��<�ɵ�\�4�Gx��|I5;Q��d`��B��R���3[9<�0����;mBav6(�� �+�V�v6�c�#L�d�qqEm>͘�R��C��)5��owN)���0�������u�AgR�퉥WW8��]U%�c�*	w2P8䄎�SO��;cp�T\Ī���*V{���Y�t��D녟^��q��{sG>x6T$DT+���/�wRܡ�۲W'�m����D7�ZK�D��z��d٠�y2������9"<��!B���aG�����KIw
Mv�C�Up~�"��$2����^��Z$(�<nGȼU��!�Qn��hc�H��B%u7[�څ+`]l����6��XT:��G,����A!��D�4�ej���B�ԋv��b�(L��̻٘�H�I�ci�����jȩ��/@��:9���kfv<��l� 5��>Nɟ����������0�a;3"�[S��aDx?tP���u�݂���.���+�FKVF\:�ݐ��P�$^�g��lcc�t���\�	�k�m���OO�r��W�K�#(�(�e�w��5������"U���Z�'`7:��A��O-�;=�� �]@i#g���yܽ��6+c��$�ν���A*?��H;y_"�V��|ê���\_߿f��/�Uv7� R�Z>��=*&6MUV�r����i��v_��=��=Sj��6�Nv���A<T.�xLa�Y9
$�,��$��z�
�	���dF&dɵYU|ße.����(��(�#�f'���ڢ����:���qI�&MQb�Q#����������[���جib�}�^` �y�Y2�.aJ��X[���\�/tK�A;����}���Ѡ޺љ&��W���Q��@���K�11���r�����K�W��� Q9f�+m�	�:��2{#_�����n�H1%n�u?3G�ƕ�3�5��i"3�G�G��\%V_=��A���R���/*pT[:�z��ly�xYOW�jﲻ��wφ�񬒕(�Q�6T�N�3��M������,��7鴢��WPgV����,�������s�\�ڕ�w?�/�oY�ǴJ/`6
��mo�>q�q���G����6i�K��l���þ���=���~9A0�������Kᡫ}�Ѯ86b�G�4ϣ�F�Xk^i1D�*X��~�����]��M`����
�(���[x�b�*�7VouB��	,��]N]����ݕ)�Ci��0`����������>=��zw{�8���)I{�צz���8��F*�����8��vZ�3؇�3A�힇��U���ސED"�+e�\@_�c�U��кՄ��$�'�9��<0{Zv�D
�EĈʧ�e�K��fs��d����z4MV��`f)���c.�:��i�:��ۯk��ylt|k���'̦K�l���:�д�4��K+O����A��lY������� ��G4���U�������6��!:���p���J
N�\^W���(p 5=0L��'����������&Q�/4x����4��$�<T���cL1�Fn�>Bn����N����w�Z�*qpי�rX�ç�8I��Wg ��ް�3�c������?H[��
��å��T޾�2hCI5��%��,�b�Քl]?�w�(�ݪ�~{N�g�iIWK�d��ӆ��^_��b�j@�����ڏU��ۦ}	YW��!�y�Z�{I��NhiZ;��ت5���I|c>ճ::Ѽ��F�h��Z~�3������L+b#?i��t��fח �G�ˣ	�J�	�B���D��A;�� b�C%����Qp#!��N�I!٤�E�x{�S��=8 M7}mͫ��Ňr��T����|1��.	�޷��`U�ũ����v��|Q�v.����Q	O��0
v�����G�-,��/�Q7�pxK3�#nע͌�V�A�-ӊ��˴������on`R
�3n�>��*l~Xi1��H�7�`*�Ӎ�r4Vt6��Lk:2�@zG3��mv��f���E�".��ʃ�'mBz�;O}�#i���f#�)���Rh��tg�]f}rQ��>_���R[���F�����A�
Z�8(����Ci	Ϳ˚:5=�ٙ~��;�g3ޕ���$�g�+(�E���ƿ#�p�#Ҳ��aY8i�����&Z�'�vt'�x,pD���*h'�L���g���,�P��r��S���kP�n\s���n9��x(�֕do:�d������RU;w�����@I��(N)	Њ�!�M5���5�#��VM����Y�l�p)����"�` �O���-����o(��ȍ���A���ٚmż��
(���<>���AI��XB�q�[V0(+
}�RaZ"&�cPӠ����L�%m���}a�j�l¬���s���9M��T����I>4����D�+-r�S��K�G�Pz���h��U��?��+m�
�"lƖ�-�3���\\ʆm����j����3q�u�=P���0FS�O��3%^\8c��eg�������y�n)~����(�F�9C�9BᏈ���Z�rS�'9_�D��$E����u-jV�	�5��o�����M$�D��^��/�cNZp�rˊ�hvG�x��YdJ3uρۘx�=d��,������hk��1���tT�:�/��0c�U�v�6ү8�v�WqUۉ��rYa (] ���matF����Pr�uM���2qQ�K� �C�Y��AZ#�K��WI���7�@n�����F��qj-7���ܝ�
x/�@��W�d��i2���{�Û��O�&�Q���6�}_����h���J�LX-Nm5�[�H��E޿0��Bk��ˇ)4�#*h�6L��Q�#��i	/�j�򱣘�/%H"+F~&P�=�dtñ���?B���G�ĢY�Փa:d<����G��/�k!��x��z�tGƥ	a=���I_��f����ϡ��EYoĦ�;O1�yc�4�N�on
� ���a!:�D:6}���P�&͎w4J�pH~���l�͝�~��)�_�Zye��u�N��\��a/�j��߭Z�m���T��VK��j�W��V��LX�)�]�䡃,
C��N�S�?�i�cÀ�XM�vM��+Y/k�K�B��k�[�^�c4�x�}���dqr@�O�Ų5����;i�!�\l*��p��~&�0�\p��'�bK��W	���E�wϵ�
��> �8��?��|����ë�>��'x���*��֒�l��^�U�Ox��H��ƣ�Ͻ��N��HA|��"��8Q��?��W%i�ω��y7��R�t`ٍ�2~M3|� lypI�l �>h
���l��n�;ղ�����CA�6�����j�9-��Ȱak��CK`�R |}�g��srSG7�S�9�x��`/k�v� c��1��?
��E��S���D�Q��b�p�r"�����q{?| _7F�m�x��%����@��a�l��pj��6�3�u��ƌL\�4��'����.zu��,"�"*Y?�ѥ?�״Z� �"L18�d����[�&��U3�խ��kց?(7Mv	A�L�Jȇ*W��zZ��W�?��k��w�§�o��eb]�.;�ŧ�#�i��Y�l�W��1�c� �s�����H�����2���B|��>�=־z��J4S�ѷrV������^��a�ߩ,N�쯋7'}*�<:w�+��Ⴅ}ˑ��`3#[�w���7�I ��A���?(��p��
g�Z>�s+	���hS�
�  >�^����ӛ�Dy��!x�,6<�o��]5�:ZU� �����
f
I&i�JJ�FP����t:y����j�F1��'>��)vL�%ma7{�|*O �m��.5T‮P�)�M?����P��g��l�6������޿g,��~���=}m�ŌxR�Mr&�a���l������̎.8��X-��$��W��k0����S��_j$�-W�\����VSt|�����O���u-��������+Wm4Xh!N=���[���o�ɀ|�=1q~l.t����s�D [P���F���K���$�T,��j�#C�DY;ޒﮇ�Yv�ۇq��Y�K[$�S�c#W�!G�0lt�=E���'?2*x8Jwh����Χ�Ǐ/�/��
i��7Q �RF�}7���
ɹ�L6���>�SyF�X��[o�-���߱)��3TW�	<'Ӗ��h�G�����iE��XB�3q˼9��p,���?�O��0�ZI'v���i�.H��PG�v��ϲ�(�t�<U��s��\�ly�sĝ�݉����ɡl
�)����B2��W�S�P&�Ap+/ɷ�(�ܰ\h��S����2�P��F���T���uD��t�ͨ�(� a��I�q��aqE��IOqm�;D�"S��S5!E�Ĺ	��:X_��X�l���:����6�th�7:�N�!s��Ê&���5��$����T�4�Y�K�U�V4c& �^��6�@A�_
Q`��xx_�H�K3&(þVӅew�4�WK_��R�K�b ȓ��y�qmeak/Ht�j����=cc�kݎ���F����Xq�u�B.�P��m�� ���`PF]R\�{�c�Xm�U������8
�{�[?�d���Q�cO����$?b�@@g͐��(��@g�Q.�O�NX�tk΃p*|C9���ge*�4�$ZA ZS�2✔Z�%�Nܮ�p(#�`jə�������I���֕M|�xܹy�v�u��=_�|T��C����E����A~��-�j�����C��z�T��t�ud6����*��+ȫ<�j�M����slxw8�n���i�`���52�Y##9X�7 ��{O2e�?�,����>�F��B�g�r�|�V��{h����e~BvP�q4�8��jDԗCّԙ��4�����uY��2��6 U�<���:-���r�h�)��;�aS��� �m�! [���G�6��u_�j��9�sfW�7���R�����?uIb�O�큁1D+�܆�Y,��cL_�vv�<��(���f"Qw͙Z&�Rpˏ��~X��R��X�fG���� �G�uW �=��,�+7L�kܢ|fVC;�f&�Cs9�g@|ؗ9���# T>,�#sŇ��S.��b]�M�6OfXbm����F->㛣ɩ�E�f��~!���dFЛM`(��VT� �w�guILۙ��8��Q���AY#ي�x�S����r�MZ���HR�����E޿U6�8��խ�<�H'^n>>+�/�Ұ��|���;[Vg��{!�b�̱��d���ƾ� �~C���,9ʅ3B���i�+��19���)Qj�MC2���`������as[j=���S·��e�<�
|������ևh-�\6����m�o v
ȚZ����M�xO%̅U4�7���82�5�)׶�)�_$�9�q�Y�A��-�u�FОRt��_�]*p�dӞ~t֬^��g�1�q�*���� xHL�P�C���^G���a�iJs��5�&$3�t�"r��o_6������2(�A�[�F�%�Z9Xj����a����f^�bo\e7b�+���:�XR��<����/F�e}pP"�`�h�A��=��Ẹj�M��m�O�"7�!dа��P&�f�h�����Bl�H�1x}��R�k�3�Kj ��:<f��@�<Bq��|:[���k��R�~bejB������h[�uV�*3�T*�	���ʵ/U$ߪ�D�7 >
���K8�����%��k�JC"{��Qpn'�ەn�Vy�� �=�)	�o*:��&,o{�B��Q����������	Y����YG7��(Ez�F���F��������������,}�)�R�3q��=����6�c���C2铱�������w-�ae�\�O7�)���ힳs���1�|�ѵ����A͚��3��C��n���K���~���J�]�a)S�֑ID���:0X�����9�V0����ЍR�>^���x-��yG�kx�):�1��5,Z��@R�`*���v㲓�	��:�qS��,B�r���"�%���a�sO1;ֱ;̎b�`a�0`��2D.E�_x8'?n�ɍ��~+o�ѫN��RA#/$�����XR����(J�z�ŋ��>���k�u�����.��hI�/N�۠��7��\`���q4u$M���n�;�å��.��֓��Ę���*�,��`Rt�gI��b׽ꔲ�$qW���Ę��^����\��?���J�N֊U$S+��*�(�uЮ;���4��S�R������\D��X;���)�L����_�g���~������(x�4H8mq����.�d��޴T���;�M p�Y!����/;�X%E0�1���#�gn����A��4����(Q�%$n������T��+	�؅�w[H%;���r}�t����������ޡlV��_�x�w\��~�vJ�PK�S=���F*~�"J]Si���]N��'�a!&�%�	>���R"�Ma��td|��+(���1[+H�@��E���[��ܧ�vs���t'����5�	M����zk�ڶ�`�@�Iˋ��8��Tad�8bܪ"~$@��P����W�o�r �X�~ڣ�e�Qѯka[�}��rTG2���@���R~�V(J�[�(2���.r��E'
^��'G"�\H������l^�U����p���MdCG�*0�p�C��G�GwYj/���W��L4ٱ���6vU|㨶�ֿ��:�K���>���U��}�E�ct�77���	��;:�7ҩ7N�u�CXz�kV�d��O�/���]�&��ga����ߗ+j�bu�_��UU��[�X��]񟊑�)5�^�~�� 0�t�ՈַY�Y�~��a����v��5$�}R��=Q@��	B�Xsys	��!�]��A?x.Q��o���~a�mbugk�e�s���Բ�a;�t�R��_�Qm8�`���ѱ S��=�Q=�}�q\��,J��p<C���������Z��W�3�9�Z��CZp�aa�}����o��O��GK�#��2a�%�sf��-Hhg�'N�4�V�1�`��C���@�F�S
��V�p(C@BV7���S���}�K&�(�
�-�Y������9E�Z'g�#����xMd��\T����h���ݦ}��s��w[GFj=-��#��c���zF*8�����q;��j�u�Tb��.���99 �����8�}c��;gxM���n��y��v@�H:S�Ql�'Z��GBH����v�M:-��������1v��)�,���B�z��2�!�R.�~�c�禙�G#�SΒV�!Hc��� a]~���r)}H7��z�Z���N3�]v�J�8�E�-e@�җ����J�$� ؅}b�����zg��dgہY�[�ץ+F߂����P�L�t�ɜ;uHa%�~��h7�裺�w�j�EPFaX�.�#
��#j�n\|"K��������b���������K���� (���FO\]ұ3�4� ߞX��dw������2rY@G6����G���ۿ��K��u��S�NbSV��R��ǟqR�\E��Ҵ��gh���	-Tc��4lt�?s�梽�ףZ��i���O3�MT<�«��w�-�({��S�A"S�(�2T?���ËG�~l�|ޠ{�I����Y���peRW�����D) �8j����(*0�B�EP#�4�Z�/�l�p�_)`VM� ���`l�"Rv,hW�eM�ɧC����VJ�|G�Z}}�B���O8�w}�E��f�GM��L�߮��cS�Q�Œv�Z��!9���q,7Z@lt~\N�l;ꇴ�S��Z�`�Շ�P�R=��;���8�U
!��N�@G�'�q��B��Yv�M�V,qrX�e�I��,=��_g�_��%_�-²"�w����w�A[`�$p�j<>d'��7Q6+�����jܣ�ރ��n3�.�A��"s��ѳwh�8�0nؽ�=V�*�?N�������U�t��ʬV���
,��O��;����n$1g�2H}�O���*`FSZ�����ĝ)�s��S��ފ��-�ýX�Ӄ���h�ǟu����Y�3��ͲL�Dt;�9��Y�� :RA]2�TJ��v�u? ����W���O��f����9?��
����?	T��@䗦 �!��a�P���y��Y:4Ӟҟ�|"���&��n�4q����tйذK�rL������n̦AT��b	0���%����M��N�i$֏�1�<m��d������p��@\�c�J�Pɳ��F�1�Ͽ������B�qE�O���!�1��6P�t6��Ǹ�
LA��I������v��������g@b.��k�2�8nc�+D]N���9HR�x*��y�S�Y�C���埮x�Ο��bĄ���cY�P1�o}�%��7�DS���x�65��a� :B_4���N.*Z.Vo�R?Ѧt�]A�z��>l��I��3��h��+N�YQ�x��wJU�ݛ2k�9ea�5�G]	 Ab��C��J�P�)%��Ϛełcׇ�'@�aR/�����6�!�?&�F)i>�$����v�ں�z�TYd��0W��xx�с��;u�'bA��i8��* 0k��xӨ��G�n��x��R�^���.c%̽������H�滗��v�F8���;�Z#O����S����#� �E
�;����C�boJ;�ķݢ[	��}񋣉3�������Z1��Py`x�@>���vߙ�r��G�h���3$��,��h��h���v��U|uxnyf� ���G���m�W���"�/��~��q�U�v��X�/���Y�ύ9v��z��9/�� �@���wuJ�"Em'd���K Y�{�|/��� �O����!��q�%.���:4����G疬'+�Z÷�H�=�e�Ď�ח>��Eut�5	���(}��_	�`�>�Uh��f�MMr���/J�,!�y.�͊��{�#�{�*U��e`}m�M�k))�4�@n�0��(��9T��}ٺ+�X�M�1_�7�:�b�桨�Є����cH]n�Y����ߥ��@	,*B9��X��}���K)�0�CFu���!F��@2���L�"�P��5�i�5�]	G���[{�h&^|��'�	��_^Pa����L�����.i>p𢍴9��1�"�� ����Nfb(�EGT.۠;�w��M�|ȳ�4aCU��!+�T56��P�ke%�������V�V�v����SB��NZ�;9n�ՐnfQ_%M�[�^.���H��=�=�����;����+) �<�_���$��bi�d͂�'d�����s���AwFaؿ�l�=�����	����*�A��G3����W~[�/T^���� �TX��6*E� %�`�y��t8<�<�Ú�>�ۜ� ݖ,�E+���=������@O'4�
#O�yz 7+k<s���R���mm��e��� Aլpo��
:�|��e4�!����Q���.��A����,�\�U��t9�t��8	����f����$Ը�q����<?-}S���M]w�T���_���X�P:l}[�ü��VL��e�%Z�EYW��
����GֿŪi�#7�B;�:G�/�i`�8��d+$ʺ����#�����r0b�cQ�6��������0��Z�=y���bR����:y����̖�ci���-�������cp��b,%\ˡ>�Ux�;���4Y�Ec�8��m:R-��i�����ߜ���J^�rds��࿯�܍��)������jy���!�"�,��
�*dN)I!��tyA3-X�����9�U�id�!��ּ�=Y��-jN�����>����Z2=`#�T g�(SR�.K<@�``u&�h#jv�n������z��,K��Uz^���}�o�f#���o����qo�C�Ia���D��Mh�Ub�S��(>,`���ө%��H��=>7<0��O��PU*���n��̀!�%s9�zw��#���*�җ6�щ����r��ף'���V���f/֐�s��S�hS��%���1�Ac:*f=��KU�E���u ��MG��(�
�?�i����!��=�S�'h\��P% �~+�o���yj-GP���n^ 2�^�r��F(%lv�7ȉ����&̾7�����q|��I��U�����N�$�W�F�j���;�f�Y<DW�S�;H���l���NQml����|��<nq����U�]��'H��?�R��Gg���ݓ矧JObM�fV�����T�咖��,�!�_�w{Eh�>��ԃ_�����$�x��Y��ױ>�/�;%���O�Ɩ���3���Nʒ��@��4 Q�H�y׬�*}��Khõ�r�M����{Q�p��9aȻ#��d��ſ��.4ʯm��_�BI�ṹ!�9@�ů�{�ڪ���А�#����8�vG��3А�f���؂�B�c�sA��vrb+ўTl	jy�,0�z%f��,<��o0�TR~1/��qɜ�N�RO���2���_E������G�,�����@��'�n�W��s��?��BV|�I��";:t:��p�Y����a

<hPo��f���67�v��)�����i�� W�2.ݵN���\��R3ͭ#��i����!(�F,';�ק.( ,L��_0^�:�PN���������V�|�88����*�ycփ� -@���, �,����@��A�"�p,c�%���B������Ѻ.	SZ��]y���w�b0����ᨚ ���:<����{_8���GB9]1�AR�w�A4���{m1�]uDt��cʫ���N�%����%���mwu4{m:�r���4�����Տ$�8��a��Ԭ{t���Qn�9%��F���)�X�N�c~���
gT�亣�DR�՟�\7P /mh/
����_��P6A����)�ձ�s��uD�G1��g�J�k�g�Y�;�r�G�7�U�����|���VN�Ti���{��� �1�#+RUЏ!U#���̋n�1���c%e�v�?�>F)��0�9Y\����\� kHL������\�v�e����M%x� Z$��75���g|��1s�!uJ�lWq���f��&%�u���f��":��y J.�(��W�!L�g����+9��2ۦ���VP�ߪ�l�w8:�{�<���eR�R�o��3~��%���P�%�Y�hıwX��盩���\ �ܻMe.�9ج�tko���E)�qbxJ�݊�+��qO��VwMb�Ư��B�J��1�b8��`#g�A�P��\9�iuF�@ɲWlŠ�`�:i������bnIE���� o+E{��.�0���8�܀Ϧ�)f^�84r��˾��@1x&��e��&�U��!�M��-�#c?��=�����~8��v�e�m�Yu��tQ ��ŷr��8��H��A��N��2kc��&�i�����CT ���r}$ϭKIwۨ�������۞\��`�H�y�Qe�I�J������cԭ�Il:����k�kCDHGu-��Q��2�>���`.���V�Q���z�݂��I�A�%F�,@{��-�s͢!�}��O�75)�qx�6�������j;�MO��F�2��P�>%�n���<��+_�p�Z��>JS��Fgd��}6�`��x�������yy�������:k�v��0(�f�����/9�8 f����+"�N�T0���@j���(�[�G��Qa���_m��@��%�K�f���R�����5����o�O�Ñ{�$�ˣ��c�S�6\�5hqv�vł�S�4�3;F�|���>��):���V��>a��#�!N�D���s��e�*�F��,���$\�Ĩ{�����l����sC�*9��Z%?�����-2wK��@oH��)��y���ň�sy�������+���R� n5J��y���ޢ���s�i�*$���+e���+��㉿u�HSX�ja��t��h��Ʌ]����1)�:�����Z����o@jܱ �<'L�Hd��� n@�Dn�5�ۋMR��u_�&`��(#Q���N��V�މ����v��lo:��%��W���B�$�e�X,q��Y�\��ܣ܊_��&�^���(��-̌�.�Fi^c�?���{~���p_s%�@�.���@�4:�)�v�G�q���{ܷ�N��{��605.ֽˆ�,�Ŧ�U���)_]��m��y�<���V�^��;˷X|`}6w�L��:YdKIۖ��]�!N&x2�ض���$9^6U��T�xOlUq��2&��_��.`l*n��`�<����L{!=�~�����Ⱥ��`1�C�Y�[Z�־�E�n��V�yx�Ք*�V�יʞe69 �'���q�fGƯ4������iY�nm����N�v�0����9͘J���f�D0�`c��W7�Ȇ.ݭ����Q�X�'
-����STR���
�=�f�	5f�b��ɷ��|`<�0�N�`����ɅSΚGTf�Ĥk���p&����Y����#R�j�"������[r:��b�и׏ӿmA�YD�wk��q!���/"�J�?��?���@$��l|&`V�zMz�׋*��p��ۢ�uį̍��Ccc��,�qg"��ߛ��5"(
�z}c�Q4�З�t4!�!�gj���0 ���^�8�X��m'C�Jɩ���M0o̐�ݓ6����2��n>�* h&8g��O��-��)��(ƀ�3�E��t�O`���w�C��<B��d�y�yH�Er	��,c�`_l<c��G�������ν2��H��os(�n$O��*}��\��WG�Hj'��)!,��~�e�k����~��N�������A�:������u	�J�is�^��h�6�{RT����c���?e���g�V	�+��˚$�C/�qP^�C?Y��fŜM�AsS)��>Bbj��!m��H>��_4n�s�#���O��`F�Y�O#���^I��ۘ���$�>k%�26�=�a�m=w޾Q�tcgEp-���yu��a�k&��136WV����M�����
���ݭnQ�-�[�E�u���Hf,��p���itBH��c&��� �TV��e���s*��T�|�������sNY�e�.C��l�����:C�/r�M�oq1kFnAω����N��,����S�h�S�I���l6X_�jh>a�|�����v0@l3A�1�8����[ 9��}\�L(��N,��$'�)7��t���3�����:�I�q�j�O(OH����� ՟�Ww;��QDX=3C�EA�D��q�ryi�He�jo��q>���@���MiNuԿ耱��л_���R�e;�6��.��h���O�Yei�m얬������j���_�����_���ik�Д���]�H�7&��c.���2�aZ&G�k�P`�k��ߺ��Ȃ\�NH�����wk���cj�藆�A��A�]�XO=����tN��W6�����-����g��Tn�,~���|*5�AM�L۹��dQ}H�+t��ǒ��L�o&U.�Gv+A��Lgm�b���@�>z�� ��Y"k	������s�# 3��2}��C�9�;�P�!�KX�MB���r�>~�
����@x&�4RW-�蛌���"�?��nJ^���j�J��­�h �$/=��Æ�ΊhC����S�(����_�_�.8k�\]��q�ز�49��Q�?�B�d�l;����_����(���H���3z�]�Oܠ_�SS�Ah��r`�U����d;�8A�Ƀq��\؅](r}5W���k��~pOt7���3(2��F���ޓ<%u�(�qo)�1z`�g����Y{��Yǀ�-�w�����lY߸�f��l��	�^Hs�P��L� ���$��²4k���̤H�J85�">��ftG�k��-��~���!���G��iZ-a����i~�	�L�������	Zx��j�Ћ<�k���g�UԱT��'gG��־�n9�qC��(������@��J���Ơ�ɢ�h�X������k����=`q�I5�R�������'�x�B��-�0� :��m��\!A-ǍY1��%,dc�O�=�z��nJM�t�]�ݲI"��L���(z����x�_j�(���R<� ��h�$�qw�HE)�z�Du���X���=���c��� ���gX$A�>�J�D3��!���7�Ix�%�O��p/��2��9��x�k-}Uc�TY��Fr_N2W-�#�"h�����ł�u���n�`|�V��7O8J��7�E���ԃ�� f^Ҽ�I�Nt�y�]f�D�H�};�EA� ��l�72�EG�U���A�q����/d�ڎ��d��s ?7�?%Fٯ'\�t�we#�ԇ�-���Ǝ.'2d�.��값��|�E�fs_=lj�m���Ҿ�B}~ J�h���\������pT/]Ʒ�V�6\	}ǯ|)i��If�[3���)1�5����@+�D�p��5�(�@�,Xm�/�?N ��H������S��`M ��y��K���=�[,$'��Wޅ
�!�g����{7	���y��r�����v+���_-�m��"�����RTM�dQ�Y�X&��ʊ��}������f����0������i;�+��5XR�>�o�q�� �-�TG���\d淿G��4��1?H0�Z�:ν���4�BlJ1����
;��u|�V���ej[,�.n�	�[��=��@4e-�yۼ�m�����JC���N���s� �����O���b��!�!('�>Z����ѐ���6ˏUg��"K�č�\6nd��L"0�Yl�&`X�͔���Bui���咏|ئh�Y4'�v"��4��]�`4G�C�Y��QO�^Ln�#Cf�w�>���k	۶&�?�>�`yL߬��Hm�ܰ�W��q���-u�Ճ�)Z�e���;
��v"���GMם��E{@^�c�Lu��� Dg�o9����9��kg��v���ڢ�w6hii{��tԿֻ;�0��3���l)	e��z*,WMIF�[��!0UL �#<����3�'b��UL(�c"�$�O(�)*�H�$����b7����-��������MA�g�Jfř���m�����-�=Ğ�{�	�I�pQ��f��NJf��9�Fضf�>��d���`'�$�r�}-"���
:6�0	�>|����|ԃA���r|��f���Kyb�ގqZ�4ar�R�%�^�V�kvۡꀚp*r�yE&���	jP�Ë϶��+�A���u�V�CY�^yFz��-�e�J��� O���KPb����H6A�V��x�]+ϡGD�
Ma�pLM]m�%��e��yX��Y-6���&t5@[���0���w,�T��vU4�c`��SP�F��e���so^�9 ���)��"T�l@�`�& &�C��5r�	������(o�|B�hH��҄�l� ��o$��ZBG�o�>5�|B"5�,~���v�P�%BW{���a"�����X˓#��
U��h(�y;�!��؊ʤzh#�p���6�X�~�x���N����;/�Z���p3w�8yi���nzHx?�M�3�2tА$Rt���hN��Q�	�5 iTNCe D[~�F̸qc�kb'=� �������s<UV���q�S��s�����!f�_4�����#h0_��[ݱ�1jLu&��ʜࢋQI�0z��}�`�a�/} y���a�E��71o:tUȁ�J�4��[�\NI0���ߐГ���=4Zy%�)4#�ry�+�o��."��=J�E������dR�䪠���2��L鋇�{ސ�&��2rU�O��7T�l\1V�Db���s��e�[m F0��I�\*��UDܸjøcE�A}QL��}����q�禹w�r;�����g֎z��Vf���s����l���Gu��̆�3s�� �4�`?Q�Щ�Qվ5#�I�WarO�QDf��Yd�ɵP�xq�kR5�k��x�>�tۛ!Ѳ���=��9���6q�wr�ZDl5!�a㦪;��BX���~S��fNq�A��˼H�x�i��nF����[c��p�����,@�Kg�(��Mf����\��;�dCM��R×���.��l����Ľg����6a8���(R���m�C�����"L(֭�������x�3_U�NmhG`�~��a>#��Y W�eH��A)�ױI% �o��&±?&��"m�SOk��^�~��f&��
 �mP�/��E�6�Z���a��}��u=�ىn�� �5σ	P����+j�<仢d΀�>؛l	�9RJ-�+�ؑ7�2�����}��K��Ԥ��rR�M�򳁧�qv�8ET��մ%﹍��i�V.�I�����O�w�t� �Q/Azhr�%~�����O42 n��Y��K⛢���%������C��_�O`��#q��Ṣ�nb���8�@;��x ����Ֆv~h��U��GBL,�1�k�X_	k��T@qd��,[ŗ��̩��h�;�.�QÝ1{��޲��\��	(d��U�����_z��E�M{�m��'�p��(%U� V&*��Ⲩ�ڐ�QY����z\td�t�·�[e��Ɇ`��`�^�]b�A� ��Ju>7Cu�P�ʑ�#�ZA�\�0�g�DS9����x����I����vDZ��������Ƴ��խ�p��*�.�1P�U��4�z_Zb�S��������9��@\}�hF).�D��|r u��H('��f|$��m�	ݜ0��x"&�p�pgTy}�\��
��+�D�wF>NEp���v������|��t�A���-���d�&[!Xy_@$�\J���)�
tV��x��op'Wف���;�LPVZ%��u���ۚ%���Z/�����Ր�/�$͜F�-䗰�ᜐ��nx1R�o���;��cC_�3�m=Iuؙ�u�}4v�0�as1z���]������|�S��d��	����٥�;��6,g!Tb�aɧ?2,�5��QpЉ78,�k��ѡ��(�O��~HB>�.����?�f�̈́����&Z^�����0�Y����&Gؕ$H��hN��h��'�y�
	_�r�u��^������t.��ͅ��آ�B�F���:,lԃC#�Ua�e`"i�� �T(9�B�P �I�Ta�?X���g���#*���/�tb%��:���O��ri��Lj�V>R"��&�ېn:�c�Z{�wAR>�V\�����r��)9�L����!.X:�0���cd��u�A�r�����20��,!�b��A���k@R�Қ} �;��;�р���542&������Z9CEA�1:�G�A�1�˨#��m� -H-���] JC�^����P������k�����(�`��	ܝ]���z����#���&i��"�~��=^J�l�3�J�kg26�v�bz��m�k�zm�󕴊:���ː�f+K���D4]�HD��=(c�!o���ؐ���A�ޠn���#K)�:W���1-"p�}�j��`d���R4
�}-��]�v�K���u����F!�q�o@���+�����g�~�S	HmC�LR(�8��������)V��?́�&�@�b�Gf�'*��.��$)e]�P˽Tr�����sHb�ƧS&-���L���F�(u� T����I�Tl��%�ӒŐ�X܋��0�⾚�b�r꺢~$^��7�L�*7�.2�K����t �*���ĺ����-��E4��CK��f��R�F�f�f3@-��+����.�"-�L�b� �F��\{CF�R�;������ǝ#a�ԯڢ4(C�°�/Ρ��F�ETX8v�m/�Qnٝ� �m��^N:4���Z��.S���J{�?�*R�4+Q�m��1F?,�DE�J($�	=���"���<Ss�E��I�YV�s��d@'Ѧ��$�R"nQ@ؽS�c
��]��E'�'V�Ly1�������F�b�l�L�Sǂ��J��_�/�n��@mM���L�@o��"�t��]a=!������q`!G}l=�z�/��gB��.�0H��֣S�r��'�T�Z��b�'%^.���^z��b�o����)�ŷ��l(��c��ImK���$�TtwZ�����aㅕ ߉��V�Ľ�1�<vp��{�I�IVo�HNNK>�-u��
��$w3~*`nN��?�T�7_h����ɞ&�����H'�b�|�v���d��rrf&_7?ZvtƼ��I?���2������S@rC'Z!~Y��p~����������t�>��X-G
�'���lМ�����6L���ڱ=H�
w1f�WsCz�ﮎ8�!������=��P*�ˀ������S��'���r��G7�}S���Iӭ���<���ˍ��ݷZD�ŉ~N�3�39��.x��BL�x��pKc������n�^�x�z�^�_7��O$�<L���� >�MX�5/��<��-�"�-|��*n�v>�R��y�o�Dc`^E�;�sE���V�>�V�]��)$p�m�/v��R4Ux����ǇF`=��#A��<���*Z
U�?�r1��cp��ܹ�ȯ
���?t�싉�妿w.���A�B/q�t?�*��q�U��\c8of���+.�$n��ԑ�R��>.����T����86�� 0�=�Z1�hA�U�nM�ե"�p�L@�� ^R>�f��0+�	�;A��PhF����m� Y�"��1�����3Q�o�>���1�ٌ9�b��jI���F�9Q3�a��ol�t����K��-����`B5Z��|1�ޱ�'d������������^C�A�:L�a/+���7Kg��M�U��m��q}�����8؇{4W�P|��|,��Y]�9{��C�C�^F��~�ږ�ь�y�&Am�gi+pe�D�	�Z�o�C:��+N��`��:�!\b��� |&*�j�\�_UW�|�@�\y���C�ڧs*������͈�.	�FE��t��|��s"�Dez�X�H���D��a� �oikN���I#�;fo��C��)�Lr�R���ŃN?�_�"F�O�"����25�o��?��)�͈]T�;_��ygv3�-�=�*�Hdx����2(�G�+�y8����:r,d<���%	D�j���:�3 ��>��O�ږ#�nB�J�s�%����"�����v�<`E�9j)�\��B�t ���TJ��K���bV��4e~қg�ϥ�y�Yt89#x�M����L��������G2��шz� �m��4��0��@�񶄇z+���f�ٚ"�I�U�����r_"1��D�e��n\l�(Ɩ����Y`C;�eݞ�F�V�mĴ��Pd(�+�H:���}R}D*7�#0�WA?�H�s�����ݘm��5r�������V�e�AQ'��'E�s�_Ȏ0��A�<�sWC�^^b9[�e�1�J�O��`ԸU�E��o���"����y?N��vɫ��b(�I�g����`��h��7d��ܚ}�́��e�Ufg����NZ�����)�|�[*�gn�&��1"�x����w��0|�˲8M�O�lU�.�.Z� {ovͷT
S��-w�Ǩw�]|�'	��Ä���1ߏ:!�w��|_)�7�p\��B}���*��P�{.�Kb��,2����l��߹M��4��γ��E�U'?m�YCk�1*�9e����ϗ�)�f<k�C����R��@��ܑ0���PN��b�8���u��H��a�N�X���3e�?�-dd�~������R�ZT;�	�y��<X@Ym�����2U!֪��|�T��|sn~?�?��J�2�Y>>5�ib'�y:�F#���0��RU�x�_��?�g���a��j�A�@B�D�oc��>J�P�k�*��!�o�a�W�Mj���ע38��3��(�D�J*�a~�]r���N.���!؏����Of��H�XCEUgq"ƂDȪu����c�頶�Y��V�]��j�r���$A�Wm�Ǯ��l���Ύp'�x�*�c܊-�lh>0�ult�4�UjT�������i#\� b~m��.\4���ĺk�/�J]�'B'"�}U0���:A��kLV�T�UJ�`�O��cSrCe�x�Y	��o���sc�'��:K�7N@�`6
C��?|L_m��;j *��U0�9tU,Yr�E�BS�_��e �{ED�� n��'�<Tc�Fv�d&�Ľ1�/ۡ�{��s1
�`�S��"��G�L���OǊ1�\��|����V��v��D����K�-��OAh	C�4w�r���7�Ht���� ���=Gp7�O�^s���:�j�w=K�&������n,h0��W�V����O%v��gf�[��FyqN�����\ ���H�f����M�Lp��e�x�����%yS�x6DL����V�!��!��[�x��!��Qvb>i�>O���z֌3��=�G^V���¶%V��d��o0g�(��ڙg��$M���.>T�{J���}��ӲS�*��&%�L�$��Z���\�uzN�����Z�� J�/�����7�����"��{��#�����O� Z�ӭ�i�\�`��?֬�t�}�xi؀z�p��uy��b�
�,4�d�dƂҤdI��diX��w�<{���Dk��yԮ��#7חT!�Bx�\���1�����N��t�:��<	�]S� �<�kˬ�*�T.^�i�4����E��u3��,,̜�#��$Wn�G��V�:�5.�~�\ݔ� ���G������3)��E���
��IY�`,��s2�+�@�c.��Y�!5�oV��č@��MC�ti�1�B�,6V(qǷ~@o<�$l���Ɨ$8H�:��c/(ɿE��ӥW�|�ס<&�����p\��mU�l@-{�/��.n��h��6#��<�&܄�E>����̣�f�Q��)/ �\j)�*�B���WgZ��8�7u6������6�t��,�[C�U��'3i�k�cߐ�#ܘ�,aѲj_]�����q����l��ۆ<S�_:1�±r�Z V�q]�	>G���[yK�8��'����L�!�P�=6S_?ׇ��
S�hI����e����Eݶ��j���SvLMH(�;-���ܣ��d��S�i�iX3��mtt>��ߗ~��0�^�L���d�:hc��˧R8�Kn�,�]���"�U�/+	��8�����V�r�	ny�\e�1m����r��m���nOhk�ԴP�sr��&�b�x� �� �bKf8��;�����,Zw8̝���iN����(�b6�O��8���I(��P�--�v�Hd��t(/�4���1,��M���:��\��e���?Db~�����"���NaB[�s D&ĚR1nN)�mU�J�o�'��"n5d�#'IN���*�P�"Q�ȱU�&  �p4T$�h'��7\�����[����QW��{Ҿͣ�n��N��"�U{hI���]A�����|�`y����,u{��o��)=P�����ԉ;�2Rl��p.��v.��ͮ��}�6շef�Qg#�b���yM���v_9>��N���3O��n@�E��Ю���b���M.V"ǽ�DHc���ƺ_`�
�%�s�=K��e��)��ߘ��q�D��k����=L!&�����}?i�PN�2����&�5�j���B)&�Ҍ��44�`B��o ���d}� }�w��H�V�a}[T�YO�.���%1Q���7�D�s2��#4�4�P(��E��m���`b����\���F��dA��jW6��ƒ�{�qE$�҈�5�vy�F4����*Ҵ2�.�toZi����o�~;��!���o��)�Uu$[�U��YL��x�P�r�`G�N������5��_�z6Uی�DY�n��}�/ R��Nה��T�G��	�2�Mk]G�\�|:���	�9������65���Xճo׈���櫑j���~DsR���Kt�w�t�����#�6�ǐN�0s��(�S������%���6�V,�{��¡1�Ws5������9�at�7ve���@�=��g�=�{�D��YHHg�B��,����TVU��5�w1�|\>��j-`oՔK;D��>f͉��ob��� թ�br��&s��>}���\���s��8��zk��+�=��A��\�*��[����=7'Ʀ;�d�#w�D2�	ή.��76!l�t�2O���������W��R���ˣ`_Dn��JU(֘J	*=�����t��	sȑ�����Bɠ>{*I��-pf�#�e��_��k��O���a
�
�F�T��Q�$��é�+�L�x���zS;�� .��0Ϻ�\�����j:�+��&}�`��G�V�ꏅ�\��ܜ����>�,ImO�H��x@Z�M��j�\������q}��Ct�@�ڊ�%�q���_���uI�����
	6'm"M��T��v�`a�3`r�z��E�y����_�L���M��k�2fI w!f�]9~��q��9��[R������δ��6v�=@��a@��g�( �����i�FtC�i�?&v�zMe'k{�7`��f4g��i�y��V�^�$���>�шN!��`C�]��d�e�IM&O5(�-9}���I`?��+u#���8��;��4����A�K��/�ƒ!����3�45l������\�>(���ri�rV+���tݬ���;o ���*�]#_tgġKI�{dPV9xa��:�/�@`2��lύ����Ѥ�f�£���X���.��`��^^���C6շ)�Z{�� �sʻ1�+hwI���w��9��� J0�(�h��6o���#�al(g�8��	H	&�)��Wy$����DѺNU����a<�J���R9O���%Nb�N��~wg؊:_���3��Φ������8D�!���9��>	�.<aVij5b�ٚO��� �j̔����w
�%q��eD;傜Y�`�m��YJ/Y���l�B�C]�٠q~)�~HT����yHl{ac�t��A��Z�f���.��������5!_���@d:�4S�Z��,ͺ4�/>�aһ���urD��:�����f��%���c8�Kܳ��;�r���D[ؘ�CX^J�͑��'e�+��E�MU ��m鬫H�L��O�W��8ޝg2Ho7���8
!] �W%芛�\:{jU{�Mb*��O�TC�*YP��Udw*fb7B��� �eCC��vw|�'{�Y�$��ؓ�C�p�y_���)��G��|�:��]�r��O��0��sǒ3�e���4��Y���[f�zW�'T|x~��x�> �����?�@��Ѵ�W+�.>�
f��t ͥ�'�� ���oYd�A�0�t~����o$��O��K�}e]/� �.9�Plj���L���\�ۣ�/�w�o�j�_5!t�#Ճ0�׌6�g��ܝ��X[P\�>l3	c���d��o�Y��+� 6/sʃ��Y� �NQy��l/H��C��LT��(��l�@[2���S4�A�@}P�i!z���X�la��'l�p=k8����m��9�]i�����O#[~\�C����s+��"9|�n_q/�G��p����tO,t0�ö�oka��< hu%�Jz ��'+������l� \O��r:m(҃o�x~c\��]{׉'��)b/ZN5��b�*1�w��,ZÓd��[4O�<M���+���!�G}�U�3��.Qh���gr��,F�=��=f��`�����*���c��d6VM��7���{cT��D�� ��Y������k}�*^�~���:�e}�ҏ���|q��~F�Ϻ��S��âb]/�޳B_ƶ��:	W.a��~��k(.�Mm��DM��p�W��{�(�^?1�(z�tD����"Ư�6�Q�wl�U$�<��½�=�F��bn��V�.1����8�p3nyW�-<�-0@q�G־��#�k��V�/�por���z�f=�s�C�?�z;��Hp'�*<�5����2��
���(�e2ܔyjsV��q�5���G:�/�{���,���'@�,���X�2���X������_���Z����
E�u��y6��:�D�*.挼�)�1w�I6�Η|AT� �̍�ʏ��u����-a�P���V�^�'�e�E�F&�m����H�#]{�ۂFiMG�@�dm6��,�s(_�ň�o	�����!Y�Ah�=e�ب'JfFhYf�'����W�M��Ѵ�����,g(�S�g>�@��e\|���&�%ڎ��>b�٣�M|��0��B٘��4��c�N�Q���cӭc����D!�?kD��@�6=r9�uf��VwG�����8�z�T�Z˝dO>vP#��.�3 �?��(u7
�D���vJ��Gr
�{�	�$��.��وs�ȷ�64Kp��9�c`+sX�OPD�p\v?9 �[�7����'knG��fL��b�76����l^�0v:s�*���}���Xa����1D���0ɺ�j�C�A:��5��Y�ɲ���?�{!�>G���>LR5:���,z�7�_�S���;�l��|hc^S�^�R���e$�:U<�įRD̜��g�����DX`�;R��a�8��>륎�V,�xo5�ߋ�k>�:�Ag��sf%Y�և��ƐV�
,�dY�j[�y��j�MVVi�S�p����.x��88��X�6RHȱ5(��T=��C%9�޲JH��HG�!��U|o
Y��H �IV���Z�Gۆ^�'k��=Rk��מ�|k��:#i��d�ՇCW<��� ��Y���P�ݴy�#�anl{f�d��*S��G���D9��=LQl��"�^S�������xf��C�c�П�e�DO�ɷ����f�&�
f��f>/:�/?�I�~Nb�e�-��/L/�Z!2���'=m�Ȋ��"Bq3�[��<�����Eyr~�{]��޺ROv�XQJ���T�����2���L�[�dʶ"�x�Y���ʅ�֋z�i�!I��#��i<�TP�~�T���>(lW�����G<ƶ�{�N���Q���9s��eoe(�p�f�6S�
�v;��򪓙���Trm��߀
�Z� K,΂B�ԥ���7o����U����T��AC��} �%hͦ�"����tE��;�uϳ)���d�£�N�\|�+�k���;/ZA���& ��6)���\\���!먶f��� �M ��VCq�
�*$�V�
=�n����fff�{�՘�Yr$�|xo��}��yn�!z�����
c6�+� җ]�ѝ��} Q��m7�����NÓ��>��K�G�Y���N�n��_��$"�����JWÎ��Pa�}a&�_��c�P��p�0���Jv�g�� L3�l=��e���$���I�HD�0����xv ��2��p$��F��"������.P�ֺ :^�^�zמ�F��.��})ۘ:�"�q���~y%�����l�"�#nۤ$�~���1B�н��(���A���W
�k���bV�ó�!B��J���=)�f����X!=lɚ�,oq��N7��N"�g���Bp�^�
-ͥ�nOYԌ"V�}��}S�����K��m�F8��q+�:Qb����c �Q�����^6
��	�?h����ש}Aѕ�t��sMp�1\���ĩ��d�����Jj�Ew*]�Uk���T���0J���T�W
؆�S^����|%X�8�ח����o��lL�o��I�$�vgn~J�K���Ɲ�zc�w��1�&h�u6����`Jib�*!x�Q��`��Ю��t�v8=<�Ǥ�6.<<[!����6ee9hp%���߄���5�Z||�.�q��3w�1
a6���$U��s�8f
��qϗk[|g��Y�z�=�ǌ_E]�~��VKݹs?���C^ӏ���wb�'�D�JZ��wos�L��p/�d؋j@�;�ީ���PZ�Qv.�~�7c� ��`Ke+����L�ۯ^� Ŧ���`kC5:���_.��}�����{���\����b/��U���KN��ƀ�;�e(Nݪͯ0S�!Z59R�L��?�p\E��`��q�P����o����8�$�hqI�1�}�߻��#�7�x>���GY(=��
sH���f��V��:��F	������}��3+��1N(�눿ta%�%^�<G �#����E��g��-��aún�wέф�}aW��5٫)qf:l��t;�և�Ƨ.��.�\��j*<h��b)���(pvx偦5��鬭��.7�����*+Ǭ]��R?��ݫaO����Y�	�e��ZHn��CqGg8�� *>-�kJ{��Z��������c�.�C�z���zJs}���`\�n���GkQ�;j�W�������\r�SB���	��7B�K�L �"D��{��NS��y�%}�I��U-?�5�G1E��{����@3����s�=���KyZȫ�b�S�lF�¥-�,��~>�$<s3BL՝�B��� �ˁ�P�MT�����uOAj��#��Z#;V@��pן�����%s��,��#Z.&���[p�н<�8��'�:���Z#���M�[�Mϯ�C*���W-����RR܅�#�v��}~�\�]�dz5��}ԀXz�u7^�SD��@��OQ_w,o?�-��pz�D�Ӕ��5w�_籡n�䅹Ϲ��9��ķ�R�p�Ƙ[1F<��A���=Ұ0���4糶-[u��b �4W�7��ɚz'GP;��|��낑��]@UӍ��a�)M�� � �p�N"_]f��t��;ϼ����*$��ִ����![x���Ͷ��1=:N
�8�����Xtr�Q���&3����M/��:y�}E�6pk�9gN8N1�b�r|��E��Rlw�aE\�Uq2u9#����"I�
�S���VƦob�����6�'�,+:��X+�5��O�D�"��́�����(TwI)C$����=������K�ؠ�����e٩k�%PG�A;d�3�@a5&]û3�C@� 0=^<\������A�>{! '�q�J� 3b��}�qA�6�]����=ȥ̮�cV%�%��Kԣ�l>���j�z�O�|��,R_���8�:q(9������ ���*xh��y����]��Ey���Z�V�Q̀���ݼd��вCc�Ϗ�@����_�i6b@	&�pԽ�w���
�Վ��%��	߾��6��d��e�����=-*������)�����{��\5����.XY�oEɞ�G���'�D�nMj��+׋2����̏+Ea�+��v�	�Q�8�Nj���c�+* �q58���H�q��OyIa��0����?���Bk	ZW��[D��p��7�ӂW��Hw�X�t�!�C��W���V�W�0���P%�$����H�D�`��Q�R*�Q�eؔ����a�T,�cG2��A�gm�+>��K��('�%YSà���4wHEBF���?�[Ή3��Ў�O�˴C#=z ��r�������0Rr@�{o-erã���z��"]\q�C�<��N�{^6�ⱹ����Yh�7$�D�"׵t��k�Ey�.�曋j���TH���Q��@��o�[�ӱZbX��{Wm��N%����2�"}6P��tH�+�t�Cp�I�Љ1FG�<�+���דh�/�b��xF�����j��a?a7��\�"_���!�:�����坳�U�Ă%���_`�d����5
�d,��U���Ŧ�h���k޲h,>��Y��
�,�h�O�OC��V���B?"������2���D}q��s=W�n��K�䲱�y&&��׉o�I\�	x ��@ ��D�a;4c�6g�jh���6L�*�����\��q�A��#pe���R�����[)���J(C@P�^e,\��+�q�m��-~z�O�!�1g�\wI:�\L�g&��ߦj������P��ii,I(�H���[;��:E��uq���3U��$���纞�j( /8�=�-�b��
�u�p�J�~M���������^�Q=�"�n��V��L**[����f%��i�r�<���c���?l�k
	����a����(k_��y��U0�����U��? �@�p+��M���|Kߦ蔎:��fUG��)�5_1BS�w'i�{s��[!j��$��<�H}߼��_��F%�:�UX��b�7n�2�a���v_��B=\%j��[�L�\9ƥ/�Ћ�khP_J�S��q&5Q�}H�R�1�v���,0\>v�!(��!�Q����XS��J�%��h����H3�6(��,73%�;�ii���s�º{�j4�]R�C���3|&�(���=
L�]��c_��v�$�S��w!۰-�h@]r�Nѿ)���R�DA��:Ԑ��D�H����k�'u�[��',v��r��G�!��<X�a<��M�֓�K��o��]x\�K5�Lp��A8���	xͅ���/�M\_��dw��h������p�+�J�t��gf�Bi�o�!� �)Y��MO�BX�]R�nf�\~V�L�H:{N��.M�[��Z�^�y̫_��V|�@_������q���W{��%�����@�bt��?Q�J��\��9km�i�|<ο�>�6	&��'N��"��kG\�����ݷ�c�eJpT�I7:�͕�e<���ڿ��1����I0
����l*ks����[{;P#��
�43fbF�dR�q�ʶE�A�yE3��jL��5���,@=�(��W�%�'��
	�2>�<�n-��2�G�r^˛���\�~�c����Q��q㜮���+�h��U^[�]^$�;Ⲫ��3�E��̘��5�S0o��;Z�r�;z;��V)P�k\�ǆ�9�?T�,9����=E8�0x���周�[W�S��|["����@�	��W1=Jo'oB�:��7^���]ࢻGX~�H�~;oU�(=��$��˸����M���K�m��H	��u+�\�����В�F<�:� @uBш�	�w%��"KeS�0o�O�b���1���Bi������bhu7�p�7.m��ʔDw�Ƙ�4[� c�}А������^
9:%o�?nN�/��,�����4��!�>K׿����=�,�7����[��؏y�6]��#°{�ƚ
��_,�J��d��~���`"���y.�{��K-d-���Pޡ.�^����$���,yy�k���N�:�G��W�����HW�k!���+�23�K,�s\��@`����=�#�*j�7��/��uc3�c+I�M�}��6]�P L[�?4�u��@.�E�J����$�������q|��b0�Q�xI���u�>���|�rIt���3��<�O�M<je�6���k��)n9\�h����x�L��#U�Z�~��ȇ�A�x��g�mR}ޫ,�צ�����)�0L'wձ��Qˎ�]Y]��2P����#�MRCvx�>�>2"?��-�D�g���^��?>j�D}�<��'�������0����\ǰ ;I��zD1_�"F�Њ	��Cg�J7J�d���[m�^��4��;��[��"v�~[�P�V�ɸw�W�İ�к#��Po�<r� �\��v�	u���_f1�G�2�j�Z�"����� �Q��2�び���)
���l��/��S��5{�DPR{2V�0� �+�KJ$�%	iƢ=L���Q��waV2�����Pl������3vp�9ʃ�m��Ώ�cA��7T�&���o�����nv�9��+�s��.��{:�c��w�4l$bW�����y�d�S�VVvn ���ow��&����`p�nwqH5��E!�����E�O�4�y�� �� ���ah�4�1��(���n��"���F(:�״�E����PT��>����R8���t�3���m�`�{L�5.��ysh�o�1$���zU��g&��PAY�M&6s�E��TտI�S����bL�s&���/i��SK����?]/+-~9&c���NzOu�b��Q��[���^*7�����Pz-���*\.��z�<���ǞK�=��Z?=�_4��t'�����<ܷq�^�^��3��_2��D�7�e@ٸ��l�*�-�|� ��������#0F�4.mH���,��CS����[.�&������_n�p	t����#�M&>�x�v9Gޗ 2
B���9�`�Wb�����
��c�e�vFb����P#=$�/����a}'>��R��&��9M����êx�AOq�H�b�z)e<*D�n�6�D@��������R�Y!Jy�Թ,Y���&ۛZ��4��>�� �3�wd*0F'��Wdh`��"���I$`�8`�`dU�B�a��r5� q��;;��M���V�G%t��Z�3�$Z9 ᠁���W\꟦ī\Y*��L3�ހ�i�!�&�Q"���uf\�ԏ�"h������q˟UG��~2���<��d�7�d��vN��x�`�)��6;@{4 ~�Zp�<�.�5i��V��x���
�������z\pUb\]�j�9�n�֤�E�A�f	��W���x�k���᫭����'!)����7��Z�"!fB/�md&��y�|8��l��8
p�k�[X
R k��]Ӎ���?	��y����'^Y11�	u��f�n@�1;���]�A��=ma	ud�;8$�^	�gE��B0g�z~ˤ��<��H0J<8o�|�e
b�?�&Ro�ߦ���E��{��@�x&ڌbT��QSO`����}���3�o�L��̿�'���E:��mkt�E�:8��-#������؉��[&��3o�8r!�~$i�~���SΕV���̵�"f;M��9����e̎`�P�mfo�68�OU"i�?f������q��"��ñ#1����ƫ���%�%��ŭ2A�U������2V��Y���x�s��]��jr��C�y��5�و��.�����N3�mH������	kb8PP�Q��ʹXA׷�
�l�%3J\�c�\j���%#�`��@+m� ����>�F�w��(����b��թ�'6��:^�xu=l�Ts!PG͞�)���).Ac��<Z�D+�Ӓ�\���=cr��nÞ�nP�cٴ{tzA���r��1$hd��J�\H��_2.���Q�o�Q�JUe��������W
K���vP-�j.#�V���t��CwijD�;��2u�\K�E����\
��JPŘZ���Î��.,�jg��K1���ց3�"HN��[9�9�V�|�Jp1�it �(����S�_�/4Yb)x?6#�ڮEc	K扡��)+��_�u���-jR��RV1�`0����L�ω�Q�J�=������������������6wD@v��G��[��S�<� ͖��E�>�D�O�P6� ���#*U0ܶJv����E?���
+ji6���C��) ] �Ћb��9
��>��z��B|?i_L�*'��X�7K�� p��D�FM��;0i��
F3���q��
���J"hJ�K2�B3b����j�ibL�d[�!�Z�	*/&����0��VWq+YaG�G�'��P��!U���2��l���ޝ��: щ��⍩���#	���̸fS4�v3�	��������MS��86�6^���pP	�Y搊nz�t}��S/{S��ӷ��Ճ�;��]r1S>����u3��Ζ�z2�8ۉ��2wd˒u����u�M!��?��b�^��5�������'TL[��y?��8rfi�2!_��sb���'�� ���3�5��އ[9= ��K�>���jGߌ�?v�5�l��T���0�GB��DFoױ�3KX��9�(�����1a�|i6/�L�����x��� ۴�ǧz|'{_�\�� �͛w����A$��G��JbS`�p��X��@ѯ��dq��Ũ�s�Vڃ=�=te���d������f]\if66��I�|n�s#��]���-�V�]ar��U��Cs��N�Q=��u������R��lQEj|~����R$om|���#��3�t��x"�o�,�Ex�������}�Ñ��vИ�l1�zǰ�����^���q�T.�ac��ѭ��rSL>�bM��t��:
����	Gg6u����,�4���Rz���l)���q\
�a?(l����k��dr�p�T�d"�����{�ǹ1��SWN�C���o_e�ה�γ��˛K�#������m.5P)�||Ǯ������|��v�L�|tbX���:���KЋ�.��Sf�����_8���虃=$%m����$�=�������L��G
�� �"U�R���R-Ϗ����F���4�]�"� nZIZ0��,}��F	�6����������xW�ż�U`�h�.�k���b�@Z}×Qi�w�Ā���/�lI��?�>��a�Lv˔�$��YV�EEZ�����j#v��ka*�p~,��c���1�[
��p+��ȶ��������߽T���|����* ������
g�M�ɨ�73�<��ӊ2�����CX�T%�]zb�C�*��,�r�/�oQ�y��-ߊ+X�E��i��U1?�@�a�@)D�2L�TT��e��}���#хt!A�DDg��)���}���l;w�,陀'ϼ(�B\���$=XkH�Ӻ�8!��͖ٝ��bW�}�6q��C\��U�Ā���Wn�Ev��$.@8��Tz3�h���辸��!���4<�^��V'	����K��(����"���R.�7zP@v���.�D�S�B^ߍ����Dbn��������^�|�A� WXer�ہv�v�##�.i{�ɗ�q�W�<���@E��Ɵ #/a�T
���&\b1\9R�=��ҍ��ҥ(䜉@�d��9km�i���*\��!�#Z�P4�A�{��f�Pç���+V��n�ȵ��ܢ�3TRK#�9c��ksz��|U9�ب�U��9O1�����@,wJ\�$�p̢�}r�{�m}����Wnɋ�`�a:���ʫ�婃k@Q\�5��xo�����&����^��qd86�B���(���L`3t��Z���E���
>>�kN;AM��u
�5��5�}]TqN:�D4���uA)!@I�˅<	a��0�֧�����p�9龉wp;��msd4Bg�d0�����[��_F-~����x&$h�r�|��9�^WR�P�S���w-�?�Ctڧto)V��
���_��E�ω���}Z�@9���z�8T��z����b���&d��~����v3��Sb݂�44���A�-��|_���B:9��M�x�3�cƫ����N��Kz����o~?�M��OP���Ht����A�mH��)��3��bK^/�����=_�'��XzK���;�򣮏U\X���`���B�� srݱ*�Ĳ1W�rtR��wC��qr�D�ۜ��S@�\yY�Tˤ��l���u��5,f�� ���o����D�a�P 0�4�r�{O_��C�>����)�z�@Z�ɞ����a�-E�{y�m�*۞�ڷ���Yv���@L��8ޢ�f_u�S����Q+�;�g씧��勉U5l�+$�̇�U�A6z�Dr�������k�z�P�5خ�X)h'T�����A�{ ����}X;��S�+F�J�ͼm��"31\[��F���LisP
�hw/ӗ���~'���D�EO����źxP�����߿&����7��ĝH�.;����o;Ԇ&m��w��1�6�«W��H�	2q~R��#�G��H���T�g��n��O�tdbJ��)�"-�i�Lޥ��TH�2EN���k������A Wvҳ�T>���27,J[� �|�e�wqŪ
`�c� ���j�`�X�+���k�+�kO� ��Nwfd��5����e�n��	AZ�!�L3�7�h��7�RB�YI<�]�x��8�����:�<�G,EE������>+��@7Q!��܇cO9�^�O�P�r���z/�K�'N�z���.l �ɫ06�]9���l�	1���{�@J1�C/uʝ�8c��H
�ש�D\|�B��c6��}�*'��ܺ�u����c��9�G8�}L��f�JVϛB���8o��`�e��s�g���C�%V��U���/�w�M���dY1ԏ�iX�O��YX��%a�����mw��cp��0g���P�P#���ue�l�h�$��Y�#�V]�B
ٽ>>49���gj�s�h�D	��`��:�+�3@(�r�%�UZ\�؝<�,o�p�r��E+H��\tQ�&����q�7�"�o��r	�i�H$��̠삾��{J����\>۶�2��Z}=	�k_�]�ĊSG�����a��o}�y��[�apU?��Ѳ)�21�3#zO�c!�<)p�`4*�_�cg�B�0u��'QU(n�_� ��ŉ���1�\  �瞓�{Bd��y�Q�� ��D��f�Z6<Q'gI���J��w�J�ި^�	vQ�v�㣠�-������8+F�10�t�EPk�^�M��ڽZ����^��_��1���z�ܜ5�KB��S�<71@��;��*�S3:H�h6��m���}z`��\q&`�>�5�X�U7�� }���1�cqm��0�mS�7�2Gn�udZ��\�nW1A`[K=��WV�3'eo�4��"�'r_�`O����	�up��<b�p�@�a��|����p�z��ĥ\�B��F���O���J�o� �xP�j�K[~�\���擾=Ӟ<`��&�`�1�B&���ˋ����O�)1sߛ���2�)��T���6L��Q��e�-�и�AG]�9�N�:Đ����n�(��+��;,�Q;J���j|�#�׾n�(m;Rˌe�-1H����J?/ˬ�h6,��<��)%vYxV�|fGG]u�h�ރ�e���i�B5gf��_�J`!ء�+"�B���X�or����Н�<�������(*e��+"�[�c~橡r�l��5(����U�U�#蚐R�S���4L+�wJ�73X�3���������.�M�g(V����ڇ`�NfTUY������j?9H�m�n{�l  `zΑ�x+J�B��G��mk�.�B1޾�?fZ��������-Rm�"��'Ne�6Ya��s{'C�����zNd��w�I��u?o<_|�w���{��]����ƥL3�]v�F`�z^��)2�hͦ��}��髚�Y �W��Ӑ<�T+z=Hc�����E1�v��O��-��c��
܎ݠ^��l!�^J���ܳޫe#"�S����<h�:-fFȟ^��
�U��=�h�5�k�����_OPl�S�,�|��-k�� {;q���������N�9�9�` 7�b2�E8��/>��>�s�6��~z��cG�j���w�%�x>����� �g~&_,O(0�?0�N�!�ODDZ���!��p���
�u�MH�ӉsUs/�� #N�m�ܤe9\i&	�� Dq.x�"m��H�Im�3�, ��i�M*e)�zu�9E�2i��OnA8�����G4$��y�8�k����g�'a�����j-	QY�fR�Gg�}v�:�(-j�~ѾK�6(D��p+���\���<fo"�b>��ļJ����?���\���ՋV���1���y�R��4h>����Cp˖��L+*��Q����~6m�AzӔ�jȉ%)�'i�-֙p$4� 4-|�k�������Z�����"aL��ݸ��lNk}��{`�����%�~�(_L*a�:7����n�V�u.:�Y^��ϳ[2��	�>p��ԙ�{��-2�/�Qڷ)������9n=ǩ�e�&�^�QC�������f�.��)�aʏ�,{[�&����U�5��n�i��u��LV׋S�6���(�wL<$���N��#I�w����an����N�!I�sL8.B��#�����b _�5���F�B�y�c,�A��P��,d�SaiN1��ʖ�L��{Rk�d= ~ F���2�Fr�P�h�+�� ^y?��>\�y��2���P�Ai0�{c�"z.�>�&p�6�K��1$����f��䣁����9��Su�
)��Y��!����֐���{�Ps��2so��K��<s����>#�D�s��&�'fA�S�}�?��Od=��0��sNW19��Q
+O̪�5�d����P݅�^�ݔ_
B�L#8;K�������ݾ��ΙO��ܡ[�E����F�fj� ��d��;2��4�<��3=�f�Z�#T���]��C���޻ \Xc��=񛊴wNz�lu�{E7�^S��D��J%�Y�<.k�=�=��{r�|H
��9���'��na�wNÄ��G �i��>q��V���j˶�멊���|�&xx����܌3[�Qm|��6�%)�{����l�2��1��k�g�"�������
�����ꈘyF��*���k[0,J6p��`�ޞ���]r#E[��s|�.���D��b��n7���8��2L�D��V��i���ϗn Ӫ&M�Tm��&��vDb����[�����jɥ|�Z>Qm�t��k�V�|jԉ�O֗Kر���:�[��mͬ	�r:�~�bܻ2e�0�1�`�x}c�o���4�&�ټ�C�Ҩ
�b�� �+�@J�P9�\���Ĥ��j�Ge rZӜT�g(,�7 �p-�+^�o��FE��2�Q��(M���PQ�S�j���A�^}���nW�z_	�9)�q{�ؿ��wچ
*?��]�X�x@����^�)6>���>�ޡ�q�a{}M�!�_L%�/�q�oG�"c }gt9��չ�|n^�=�p��h<��Z��)��c=�G4��ri�q!f3�'_��E]��Ϯ#�gG�����r����s�<Z'��ŗ��~)�R�:c��5��s�l<�#Xq���Oj�j��2�H'N�1`P�B�W{=?�
}�!�� ɤ�>cs��kλ㶲x��pe�âq��+<���U͆ڇ�F
jbm���j�Ϟ��4��N>f9��$�q�%f-�R^�6�^��|�!�\,d�C ^�-k�O��
�弌��9���'zI�0id�^?*�%��0@�L�a��K����H��/�U<V�F'��!�^7�x�"ش�l.5\b6��z�*�O�O��G��z��A����c���]�[�Վ����)�X�)����Q�N ��H�-�`�R�U��k��B��1E��.�ONV����8!$�y9�k��:��?���G�r9���d��.�F���lW�XĬI�걛������l�p����'C�qz��x)}�z���~e�ҘAOa�%�<�`$a�^�BN�P��p8�����!�Red:P�]������1&���`�&����2��'6�J�Ǿ�5$�gFe1.6��봄���S��K���A�&��d�EԐ�eɛc��}�\s;�
�%{�J�������l��7�@��g��AA`b��I0}Wto�,7�>M��R~�����G��G�寑+]��u��.l���Ң��������8��o���|3��5Z�|83`�#�����l�R3 ��d���S|d��W�F�Y��~a��ɜ�z�-�]x�*#�T���G� ��.����L~)�M�R$��7V{L�$�����f�p&r+�L�/���a�Ŵ���Ke�g�+C�TТ�KU�D��{?ҿp��32����]ʖBY��	ϗP��T�n�r�*� `�zm�V��H�'	���Q���PBZy����
�D?�9}�b!�����B�(�i��~�! fŝ�ջ�r��ߌ/9T2�tK�<ҩn�d��c��Fr,�^�#�P.wf��y�jӃ��'����饱�W�.��>�S��h���F����lBՎA����K-2����T����M]-��W�r_ýʩYA�H�(�i4Kc�ă���g:n��΍��MC���(�춳H0&����D��!d���ݚ/8����	�H���.�Y�4��qA�]T��d'_Q�����ĩdZ�M��Pe��-,����S��p�Ra�T=��^�xb�#�/t�=4z��]���7e���}�B��ԁ�%��ly���:r�'X@v��Ui��ڧ��x��v�:y|�{�_�Pל }�)����?�y��iT�έS�^���K��7�TZ����Pvݭ5���8Jfa�e/���F�BCM���Q���:(��[�Q�@O�W�MW_d��!Mc[[2ط.�����K�b��{�G�0��Ճa��c
V��A��Z���C ��[��`�����zN[���tm����nX�u�BG�]���$��I!�J+�b�ڗ5�I'	W���yf�_T�T�C�� -��6�N#)�$��s�n�+��_X�]�'��Do{<i�f&���h2��5>�� _�˙ld�4�B=h4�v���fVb\a�����`T�3��q�q�����+�V��ST�E[����&�U�P�s���o�hn�nגF�7�����ozG��y1:�L��rKɹ]���F�w1&d�]�6ժt"��Y��I��r_��*�D��n�`FDgi�]���44���C�8��{�S�W���y��MN�%��P�KB�1V��"=���:�_�QŏO�? vݐIr��7��@��aq����0���N䦛 �[�lPR�QW�JEIL�y���NH����=F�O�tL����j����� {ǂ�yي'�����_`��‗Fd�����)�����;�D�蕯u��
є�������o����Tcx	�/�^���<p�/G%:�ul����mgeYe+���V>����J�9>$�̈}���l�E��	�h�����x�M+{��[�g~z%r!���6:)���/D_��ٔ��;V�L_6@��Q�i�R�
NxQ�����w�'BX�u��I�+�8*\��6�:/)�o��hѓ0K�,���E��Vn_��L�NT�
Z��6�8Y����R\��CL�j�ܲ�R�-�r�>F�����M�RIzԙPk1_E��hu��v=!�B~<���g�5؆�8����W�Ҩ���Z	�L* �Wb�Wۻ+��r����]�h��|�X+�Sh�YzoYD8q��g ��r�{�uI�v{���.��洗��_��&\5���i'B�G�73K�K�+f���{�o=��0�)���z������)B�=V��+8�ͯd����нl?�����;��{6����t'�����9h;��?��(�)C���,��5�� 2`��������A|h"�rkN=a���]Ժ�j���W;�Wղ;p+9��Y�$"��W��h8j"j+�\]d%f��x�����\/7�lU�uj�*[��oZ\�+���98��X�ܭ�D���r+�a�ӹ���k��y��#�l����I))���l��ɵ����]�_},������Z��VԼ��h��I�KR ��6��殀D�_�尮��&�_��uK�;��������X��h1xmm)�J����ˑ��lX��d*�V}��U2q�B?t��'_7�KzKO��3e����d߃����FO],7�6�r�u`�+�v�ݔO����ST8/���J	��)}����5ݜ�.����u��G'���W~�p���1��cEEoaK��R��]�*�	���|�,;��F�]�$�s�Q�kOnö�M��M^�M�a�Ec]�����g`e0Q��o�|�-�'���|�#-�+m�ZI�2�i�ؘ��Q�"�e�P�>b��� ����8���M���?E�.�wak����C@|��M����yȻ�7�)
dn�N�ѓ��U���W�un/��OJ�)pRș����B�X��x��Ku�ϲ����IJs�`X�ks�(Z�V;�ƛ�7ga�&rb�F���2~z���|���S�!�����Ύ�Dg��`�:Ƃʝ�O�ËS?��

�w�����Ɣ`
ۭ�nH���S��E(Q �=���j�3���̀QgÎ3�����ыV��I~.����
��E�	\���)�_$F���I�&l�Y��H�hS�-6��p�JX���4Cwu���1%C�9[��������qu�1��4��y��`���]KO����v���Q�V���M\�t�T�U�a|��U�}�=hM�2�0R0-�^����Mu���x��Y���� $/������4�05rC|�"7�^VBf�v��MUֿ��.�7	�L&&�x��ґD�����u.�av�/��i�-���|4(W��b�[�N�;�����M�j�� �O�r� g	먌a$�)2 .}�0*K�Yg���6I�=�%Cޚ�
��܋4�bsU�'"�%
��J��U�įW�+�',y����?Qj�� ����%�q�����b��hX�`�¿"|�����bc>r\���;��6� S�v%ݬ�=�"�/,��)�L[�t)\���x���_ϗ������L�FƑ�h����Z��_�b� �2�5)�a�2�Nn6�l�?��c%�U�g��آda�6)�w�ٌ&���,��Qf�Ԝ����(H��u����l���P.woBzk�r��ؘ��{�l(+?II:���DTh�д그Tθ�J=%>c~W����]|	����>2E�XV��!��+H#�}�8�_D�ɽ��M��f� SBe]��aR�
���!w�3}�CO��W'ގ��2������b��Tw�C��6"݇~�>,j����� =I�(N��9�MP<�����rW��	Μ1�B����Qe�r/��l2�Y˂����B[���Ed�a)d�
�����6�6#���K��n���]K��,���Ղ#hEU��,S	ft�*n�u��ީ{	Pkx4�i7*�(�E�4u���%@s^6'&&�$ەt!�,\���`c�D���D�]7u.�8�p���i�W��~Qb�B�U��)�F#ɩ�Bs�_h�k?�bV�J�Q���5�zN�b�� PGk��o�J�>��fr>|���$t2oHe���(��yKQ���,�Nf,t���瑁kӞ��Kբ���jz�2k����V#�:�/�4���CT���'��M�������d�v�����5�e%�בb?P�J^��A#b��^y%H��'�wr^����NbߜE�����`՛BWݰ�܏�
F3���~9v\��9/zb�>DN,��1%WPp�o/ǁ�4��
��Z�VN��Ɇm�(rl�z����������6/�Cxz��_��'��������̃ 1/,�H(L�ˏFZ�h�m�������%ȧ���9��6q�;zN��AG�:�k�}) M`��%ξ5���*,�����>�p�ݗt_�ds��*�&�5_Qe.������ h_[;�^^��ô!�����^�H���͡Z�5�+k��P�F+xۃ9��-d>q�
�%���1�b����xћ�A���O�:��0�������_8����$�K�ĵ%�;T��,y-�G���ߚ-E�i�Ͼ�L� m9������_�q {Ir�QX�@�o���@d��b�;D=���"��D>����]B��FK:B]��9�I�gU�F�O/<0�h�Pl]���Y��RYq��c�]{Mu��3�B�|t�相g	��&I��6��Qh�*_|2��gp��q�G3�S8����*�(.`!���P��5cH�r�ۑ�R_���"�q�U� �	{���X��QN�m�v�cf����
��\���O�F�@�B&�[���*8\�yvaQa<�D��j�q�U��cQOF���{\.��[ȣm��R����w
�F$;���Rӓ6.�������b>���s��{��q��YX���7l�<��J���5ĸ�_SF�7��/!R���vu�-K�";-��@����h�-!��R(�ς��Ja�GF>"W����i}Y�UI�3ճ���W�63��0���VU�}��@�!iْ�914f;�׭8uX�L5P��G�_~B堞P�O�Q/���)�ְ��#z}�q�ӥ����)�жKU�46�~B(�!OʝCe�&���&�Q��GaD����3/F�ඖG4�7�g��U,��W{�j�0�YX��Z��x�_��'f���wŚVM���K��$�G9!�K�>�@�`w?��~#׳cH�����ՠ�����k�c�bX53������R�'9C���&V���O��Hb6��T�Pp�)�en�'E+%IW�I���3��:��~<��l�_.�y�u�dYߤ	i>�ΐ��D�PT#����|�)ظ琹Mͤ��(W���	��Ĕ����{��.�o�d /l��5����;���!>��"���Tx/S�fDˑ�;���3�#.���QR��]>K�f$ļ����:	s֡�����)��	x�crK`H�ٚ�/�e���=�ňͭ6�Ë��@T3�'��aH�9���L�៽�^\�Ci�v*����
�A�f8 r7zu2�����4��n��
�>�mq��%���f��٤٫U?����}���jA45��Mp�O�]�m���ґ$+���vf��@�$���uR�C�����n|1�z�5��{��&��^6����K	�IZ�,�2���_�٩�7�a�D��[䓙�T��u�7>Θǚ�&�8Ɨh�Nb(�Ln�%���9�bo�/�h�ѝ�[��e&����j�6�70QZ��=_�%�+�����QbZu�6\Hǒ�����1~�����`��2�8��"h8b/<�R��b}��Ѣ�����3����K�k]�G\Q2I<���#V�f�t��b���C�:��ڶ�^��ܐ%�s�6O3m��M�Avo��@�s
Sj�J��ӷ<��葰:\�[�V�	�7�^̿.����)�W�c�5 	֌��bG�(��mx_��V��'?�o�ޥl�����Eó�s��F������ig5'�Q��?L=�#/�p��wu�U8�u >�1@"�h��ɽ)BaE�%0�Y�*L4��0;�A�o��7u�� �מ�rT]@$�Β�>@��@�qe$���4��z���%̟��C�֠`��H� Er�h��L��T�x�}�:�}@�eF!��[��������Fm^�f��"�Z��\��w��гM�i�H���� ���th�ݬU��f��ZcC8fKq�G��k�ן<5���3
b� ��!���Tm9��έ��u/V <_��#@5B�*8��:%-�sL�����BC#=�@˾ �wFR��|�: 6'�>9������i�W����)��*���8�G�뵽)�"u�	�Y�܁#��g����p������o���� Q���[c%�~�;�(��JJm��P���"s�8�S3!�J���V�5�����GrI����ߒz�kwߔ�"m���Z��)F�O�i��mM��P��}7U��7:��	��-t��9��-�.�o�/�F��o�p��SӔs�˦rZ..�]w{�*����)(����{�_�����\���˥�xO7�K�]����K�԰_�� (E��\�3Q�=��@��_.�9&��w����2�O�d ������L�:d�|1�K��d�q�k��w��X��� ��I0��*"ɐ���
|'���)g����8���cT�l��l��l�����-K��G��܀q�_xC�&�@:�߾oJb�c߀@�IJ]���Bٝb��������&���1�����l����OQ�t��3F��V��njkh%�[���UԀFV
��f���
�pRM8]D69f���k�����v�,��n0o)D*����k��p��n,�t�ḝ�T-Tdl��DB�<�]�ưo�L:�]A��E�|�|R�~����h.=��*_vP����7Iu�"�*���o�x��C����T�/k�?�z1�6H�lP99#f��Y�Kѳnv�O��� ~	�*�9�:m��k�x|��2�?��-��E;�\��aOWn���茶�2�'�K'#L��@��[�Xwwxܶd�.1LH�.k+��ݺ�b����2J����;H��$��������c4 ���`�e�L�Q{�Ȯt�ҁG0 9|�ŭ��Wյ1k}j��xI�(�W�#��V)�qr`/�#
ޛ�[DO<խ���%"�8Ǆ�:�~�W#j�ҫ�k}J�c�?���!c˩��`��	��6�Q <dI�U���xu�C��i\�b�TS4w4%[k�z2&�$���l�H���Ft�����?���N{5�X�&Q��B;�ƽ:��Ӝ�Ɓ��@g��j�ȵ�c����r��ހ� �<m��]<���PJ�l�'��Յ_ONlz~�$r��\�B��5�h���}feࠐ"m�)�4!:V��wC�8U�I;/>�ڢ:Hc��� ~Zh��Q�x��^��)TJV�բ����붖���_ Rc�	iAԅ��>m�7N4����]�p��k�����,g��ӯ���{�]7�.���<5����x�ܲ���뵧|�7��Zuc�|�*�O���K��gfa%���L|k�$O����X�`����Ժ����}�~)mI�����`=v� �t�J㞙�~��|���ok'@��H�Xv�އ����ºB����-6i�v�����0�E�{�P�r�^� 0�������#����ݢG|��)R�2^�M���p�Iv#$�~�͚hr��9�z��%��: L��FR�H�u��
<���R��]RM���3����g6`��7�}�sT�_�Ps��{nn��� ����J��t\�!/�!�������1�Q�3��P�o����R���4��'�=A@�Ю�đ����Y�܎�j;�n�l��B����O����EED���#6�ф�f,#n�9���n��1�.����5�{SEٱd��ױ(7�b~1l��0��4�/��q=q̞[-�X/WW���ʫ����̼ՏR��2���LP��_i$S!�=��&����%�?8s𸟃�|�<2���8�O�X������s�m�?�S	�[i�7���YQ�; 
�5{7�ޥ�'s�+���ݩ�[9�a���:M'z��1�_޸��{�~L�'�I�����sQ�,�Ɣ�`�=S�5�p�dua�1�/Y�Wݫ//��{��j���YU�)k����#z��4�A-Kaǆ��������~��՘�
A�@'�^3���&Ӛ}A�0��}L�[&�}�(���a��$j.�hb��r�f�a�hj��2��"2���\����(n�܎l�]">H륞��O����̈=A5�����Gg��\���e�, �����,�ݔ	����Ff7�߶g`޴g�o�!g��������Xh�+,	����c!>���s���ڴ�H%�)�xG=|[c��F��0fZ��p�Rӿ����wv�Gm[�5���i2;�$@.�G(� ���h'K�������<����v"��vn�+}[�e'	�)om�u�Q*>M��/yvT{��֮����7�FCiH�r�N����3�"�g}�"fi��Q���2�˻F�������j�}>~��ّ�4M.B�������~3_��z�M�N��oC�i|g\�	l���l�I�N���E�(e��;� ��e�(����xy�����[B�m���~���T�������~��r=4J�$�cV�z����{��oJ̬.�i�v��N�ݞ�,���g�ɴ�d�E��J�Q1~�q.9����y=���h�F���QDC����"��bm�`k d�<-��v�|u!���m#AH�U����gͼ��h[���Ǽք���/L�]����f&,��p���w���`����@V�&�69���7���Ձ����̻��S��쨾Y�L�dSX+�b��s���E��U���5�RW�0�f�;dC�zU{�� ���H����4XC�7NI�"ܟ-X��X��wM���Ze���Ӯ���>AL�}���5D���<PY��;�|Z�A�Ib�6!�
mY���p>U��8��3�<XYջu�W#:�逾�
/�wb@�wP�J�XH�^�'�ɏZ-kN��H�ڶ(9���#CK�z��I��	��r_i�YL�I��(��T4	����S�X�"��i���"t��`
����m�_%�9��ByzյV��4?�����`k7�v�u?��}�����(E��R��2��:q��-�O�͹��I�_�9�3X*�Ο܇��Z�?i�lL��=�d%�Nq�u�w)2��^@�g��_�lx��(��)@����t����j��L�|C>K -*��z��K��k�4B6Lߓ�۬�1����h� �����{lo^~� �D�W]E7���'���qh�㲝�q���0��\īs�M<�N��&%�7�	�	U�t�H�#]ne�}EW�JK�����NN��:B����X�+
� T�!������}h���s��_��ria�=���1��*`�\�^��X2[`	�)�M��j\��'Ř��������p"SkP��<�+2MR[CJ,ƪo�Ӭ<CΈmGJ��C�D]���u|�i8�-�P�{B�M%�〲�6�{�n�S�j���I[ip�,�7���3��n�S���A_��x�oďQ.�&aa*8§��1��o�~�!=�_���9��T�$ņޖF��kI��2�C�v���o���X
�5)=���W�7���lB��ٖ�ԑ�B���?1�.uf%��U�rk�l�5���d7�c�q�s�+�Z�k�c,b�{�l6GŁ%�������[K�H��@&�+l�  �>��oTtbC1�f���'ɾ R?d�7��쮮OE�p����`�U�)�?��|4Z�h�/�۔���_Ǡ(t|u��4������(� �]��f9��+Ǝ�K�;l�	/Uu��07lE�c3�
�g����[���BQ�y�������{��p�8׋.�b�A�m�Z%�Y;�V��7��ښH��{�SgA)��п�_���W*��k3�9����}R��e���z����s=�-͖t}�sMT� ����u�t��.���U��~�� �|3E�%�V+ ����ޯ���@��cT�L�b��4fa��,Zp��{���~�!��P ��5������dz�Qv�:F�?� ��2Z��vF�Zd�4!q��@�c�Ob2�_�;�\r�و!*�0"����h���ڊ���U��egC�֑����8���<�{4heܐڇ�PZ�[�(�;�G`!1��cոJ�K:�r=@4~���C����T�/&�;W����"�~���׽�Rv��5�%�����-�A�3�'!y�?���S}�C6V���o{ї���z0���wxq)���f
���VS5y�"��c��7���cm���A��꥔���"Im6�u��e�d��	곳(坲;ڼ)0E�&��_�V�䳎�G�d�#��e(?Q3�<���^�m�#I��/Z_���|���ȟk����5��l&d_�����8�u���;cDS7��t˷kio�f�5;�
�(`)�~�|��Hn�˧�S�Kng>����kQ)|J|8���IB���v�&�FSv�VK�7@K�/�<q]aG�	 �3�q��$�"��mm6Y/�EB*��	�V�E8�Bd!��Yɻ��$@������Y�3�1~!�>%)D
��ϊZ�}��L��!�<�2A���77�q��J��Ո�����\b-���yD��PK�FPjqfO�s��E�k����A�8�u��n�(0���D� ��̗51
i�#��q�S�v-0��oI�~�׍^Ra�����}�YA����i���e,P
���<@E	���T�
���l��+��ɉ������K��21W��ԩ���I��m�{@��$,���v����GS�tݛ7'�oW�6�L�Sj&��G����5�*���'҇_�N�L����:oRf�b�Z!	���me�f�AF&Xi��A!,�A��j�0P�įk"�'�.x��J~��F��n�H�XF$�� �IY:�V����pȩ7A8F1ġ�^Īo&��h���/Xie�ba`(�Hgo�pc�0�>{t�j	����d��6j#a���ߓ�.�'3�I����gw�o�4R
�K>g�C�(,-$�Qp?�[jm�~�yN��	:Q8:
��%l�ܐ�ם39����Ϋ�Ȯ��X�IJ�Y�| ��J���Y�4��sƃ�]��0[�W�N?�*'��z�=��
��p��Es�(!� �f)�U��Vł����w�p���1��c�d�O��P;�q?@־��X���n%Q�B��bz�Cg�������i��P4���T�3BNa@��L����2��`{�nJ�1���/�����sr��rV���-����׷����u��z���Xy]��͹�]68b�c��ɌE,�1Ċ{�T{[y�S��3!u�����On��h��7������î�iv��'S�렵3]aZϮs�T8E�ϩek�B��}�S�`������
�6�h{@8��u�TIX����+��ҹ�s�ж_�r@������Ͱ�L��
5�B�J���!m*w�{�>G
W���y��I�-���*���CA�8v#�#�����1E"��3�'W�&+a�jzJC^��=T4+�%.z�F5�_W����2����`B�u�����ˈ7���ºj	���R�2�Y��
��4R����|#�~�Mro�����Lc=u)�S�M^*�4�(��`;u�Ƚ��Rϕ>2)/zNK���e���QP�-�C7V�͐Y(��A�י�u��F�t`G�eK!���_gh�YU�.�wQ���Dz -q�@�N��5��nL�!��~��}D\~<:0����bb<ۻx���@Ko���Hv�w��Y�f�\���
[�!��ds�9����V����&�U���j����?�zU�aE���p��3x�W��M�H "t�(�m���{���Q^[2NWr.A�%��=_h��|�� ߀�`Ŕ\�����d���n�c��@�,2oB���\v���HWE���a���LM��X1��e����Y��.�+��J���=S����+1�7�z��r�䖱�e���!��5��ה����C������b���%	버L��8!��`j:���q�O�"�|��:�����P���<��_�L�v́ƠԄ �!N��5�KO�~᛺�3^\!�Y��2�X?ȵ�,�y��|������$s�8�Mkt�t�aҦ��K��5�ϡ&
a|�EU�8 ��W凾���4(�^�c��� I�?q8�Z�!�/�"����Q�1�X9dE`��E}���[��9ȏ����q�~O�-?s;��)8�{Nf�����,�"��h�F�5$��O�g�׏�W���)�f����a���>2T��m�V+ϧo/��o���#���:�&+��^�!���J���փB`�ñ&%��'�̢�e@������^�o�w:E����9�1�i�Q��������Z����?���
�����R)�3�s_3S���.����͏
D�ۅ�$��$�˶~C��J�/+�Ub�備.�j���ı)����b���-h�ŵ�Ԯ��R��U����vN��=�
8M�V���Υ��6���$
_.ia�w5y]�F��4*�2� ,اOu�E�V����5�	N �),ɱNje��u!G#Ȗ��5�'7��}$�I��:C�r�/�kH���3u���LD�AhͣcrZ��.U*q�5w�&�*������2Sq�����~c���$g�?>/i�G���C����M���`��\�k���Al�[��!N���"��~��15<V�7(�~ωK�D���-��I�m}
Ϫ)@�E���}BJ_�AI�?	��?�Ć�)(.2��Eʋzr�I�&%F�������y�5�Iɟ����k�X~��N�?;��rJCV<�DG哢p�m��(��12w\��<�2�;��{lX�1<���V>�B��v��@n���+�\���I�n�m���a��ӱ�䲪 �!�:�fW�i�C�տ������PC�4c&^�@�9 ����ǰf��+3��Rr5[��J=ʄ��:�}�lV���ݣ�!/��\��zA�D�Z��zƩk`�k7�t��U� -v�P�WX
__9��"Dse�4gDa=��xw㇩d?ԖR�]���ZU��&=+Z��ud�z.��Hrk6il���7��^��<�V @��ݘ�:�?F�ؖy�
�3,��E��˶��әr��ڢ���'�o���te����ȍ��ZM�R�����+~m�GI���S�.p2�o���[��� ��ʷC�����.	`��p���s�	�>P����}��i��@~����]��.K���C��0�k��1N�ƚ��5�Y�/� E�Y��$ٗG�N�'ԫ���쒵�vq���l�X�9��Zۯ��%����ʵ�qE����&��̮���<��Ԍ���My�N`5}�>�eޝ�AO��:�&�=��9�4wxtW�j�]:��^�����Ʃ31,����f
W�kn�� a"(��1Q*t�ƹ��6��76��w�)�^��B:J�d�fX�K��,���<�����䱒�/�l��[���3��}��$H%�-������`15�o6]��S��b.�s��s�����.nbDd-_4��M��]�x�쫈�U�\�&*/1_�`)�{�Z����b��p\@ov ��d��\
ń�F;/ǃ�cF*\u�.�'S�c_���NI]��آ5��X�	Z�;>=�=�H���gm��I���-u���������W���4;�9B��.���X���U��wþ��c�[�-����]
�
�&FWoW[4���u��q
���<�N.�R�.�qy�����)b�0���Kԙ�8��0��I��B������2�9<ІTy��!	�z� ���BL�@��HWվv)q��;1�g�>���T�� ��&pEz�۸,�o�7�N��,���I>F���:�ڰT&F׺o�H���֪"�=���<l������*8� ��0d_�x��_hW�W�����k�����:�J���%�9�QAL����UK�PmƄ1�xZ�B1���J�)4��RAM��k��m��9y�����2����#�w
������<��Zw�T�/��G'g���7�R&$`��h-�ͬ�U|)�n�l.�?A���!X��@`��|Έ��߯��nw�B2>�n�bj�e�;k�ҏ�_#t�����X��r�&���|���7�G���lwv�`�ut�ۚ��^������`ҧ��'��]'�P񑡅2���҄<&+��V�KaF���Uk���"��12uӭ�c�WN%�f�g���Km�P<$���9L��K��Te��$&mBe��z\tuHXj$d��0'��#X�"���}�fZ�����ʽE�iUE��)����:+��bX�w�ӧl=o����ݬ���{�Y�U:P�mt�+��Bfbc�N�+�o�s�f)K��F~��G����[2N�~kGNqM�|N��@�n�����J
�+�
����b'�bV��ޮ���JJ�mp�P�<l��W�~�y1�`٘D`���~��)�PT�!i%�ȇ6K���7��Њ�*y�sJ "|I���/y�&TL=�=>Zϩ��� ڟľ�'Vl���R�yT�j�C�{���㷡LϦ��V���I���m�jjҌu~/��{T1k1�XU$�+!�^Z�NáQ�ۚ?���:�� �&�h�d�rO9���Ư�&�>�7�'\�s뎛��SN}ځ|�9l�8��{7#g;��K!�����<fGջ�?'T~c�L���S��/���-�.��=�;��#�x�k��+gX��E�#��o2���yd����K9*��|>�V�1�1ʘ!ɛ
h�>�x'Y,#�M;����P��HvoB����,J�ݶ爉��iX�P�A���e����k�!yU��p-��k�y?oW E?0���-�T��?q@�qC�#��}҄����2��׀��K^��5*Z
Lf��&��'z~�F����x-��^��%�bfI��uۭ�N�FSu9)l6�樓��Mo��Ӵy$�<�؍U�ٮE�}�QI�H�?�L#��2O ��^�e���r���G��l�Ĉ�z[0Oj�-�oS�)�sͶ�e���3�N���=�����e}��}�"�D��-�U�0��ӴZOsa�b�L�ZQ��6��![l@G<+����5�d{�G8+��T��` �VD6�Lc0`/�7R|��`�,�I'���Ve�iM�b���=����x�*���)T����8�";}H�.8�U�W��^7�5kB�W�x��(��a�%��E��D>XO�DPN�C��`��VB=?[���潞�,�Os��o�I5\E�k�	�����>��I_�d$�%:����:��,��~�(Uu2��������B@0DaO}��u��j+��xB�M�ǀ8��O���3�\!վc�)�<N��1}�4�m7��"A�^����Y�P�5�?<��6��I�9V��*C��50��3D˺M)��:�TmcN�>$}�,�v\3�r�QpB*�AR��F��z��aS�r�X�G!43�쉬1���J�����_:��R�|�&j�n��$G�0�mn
wC�[����B;tB>N���F|�u�E7�u)ш�C�.�9)����Pk�M�l_��r����S���V�I{�NE��_�f\�j���&�Y�^eB�|]�l0v��[w���l���$[E
�Ҳ);�Q'"�~�N�e��)"�"F�|���ڪz�*.Ny���B�$��?�A���`�	�		���-�Z�h"�����'f���Ͱ���<�V>��?��7��;�C�'_�OJ� ��}�\��7��$z�W9�6�M�N�}�������2�ч�\A`a��fa��a�M����3�
�(�'�ymnp�X���ν��H��;k�m�$5�~�����RN��	7I~&� @� ��23�?�g�2i�����N����m����s^9�M�#�5��5����m}o���ZA2°�c^Ҟ��'pw*a~���+*9ғ�w�z^z�NF]�����rOx,��,da�i[�v�A3�8M�bFE.�<�D�]�QV�):��h��W*�x�\L�ǫ��1���{�φ|i��G�&~(���"9���ᆿ�b.��RX���8_����e/��|��"��E)�Iy�m�Ĭ�N�������*�-U�?��}m�D	���
�	�P/!z֐ݴi�^�.#3�(S��i���:�6�Ju�0_F���:�$\U��ȶ!|�4"���B�0��c��q��qKږ}�Wz��@��hO�ޕm�	4�I��ˌI���ɱ��2\W����<����{����N'yp�4}2���L���bo4p	 �*1S9�_YAWT�v�1�Ƌ�8���(�I����Z�U2"�[a�+�t�+��x
�9e,i3�Q-:�a܍'1�BM��d|=(ײ��d�6W�>��.v��s���N���kjّ�!�0[��;��K��yCv���r��_+��f���K���)² "�<����iIƷ�^U~�	%H:	禉�Q@Y�������^�����B�Gٞ-[�U��Y�nO8\u�Z��L!�$�Ő��UƧ������2$���8_���Z!�뱕��1h��B��g�|hp�ތ�}�R�z|Q�H�xN�^�w�,�=�o|���1Z}�#΄h��yt�����&���T&�����Gi��Dhn�E[�bk��R� ��I�h��hDB�yp3V�h6�M�����5\3'�[�@�a�<��mQ_/;���@�2�G�\���W���5ͻH�0�����HK�ӊGQ麿.�*jw�)U���6YyET�JT.�C�Cb.Ե�%r݁�2^qľ�8����]S��)nT����O�^iK [�S��a�	D�m׆��CON$�����������$��J�c��?�a;��L��u�`�FW����TR��i�i��=��#ȸ���:�!�Nf�2<���(�����^9Y0��1$�2�>�=gC}s�}찞���3�W��[�/� ����=X�\M믱$�'�jX�?'n�c��1`���c*���2ڌc�5�$��K٤�K����������'��e7��hX�q�L�W!����?C��?f)�(}��6g��b�X��#���G��
�*M?���c;4�&ڭ <g��}Wo�D�0�d�x�����-B^�:K��P�j��5ɨ�� ��(�p�����G��!�B���<1��b��^��#ёH1_�Z�c��|6/�$���lm4�Ӫ�&zJ��	�2\M�2Q�Wũ�����R��S'|���+8��n}
��^�5��)�����%ў�ʪx�*Ru�Hn���j�p1��4�S ӘmX�U�6.h�4��J�d��B�|5�>��W�7M��:��Ѥ�s,�ieF�k%?	��@[���@�3&��:!gy��Y�{�R�3(�y��e�mg2��3�B_��5�E'�`lt�M�3.�]�YT�����-*>�"KX�y�t��?ЕZ�k�p,���Gl2/�r���$;vX���Im�ʆ�1�Ќ��TG�r%G�a�|�1х�b�X��DKONTu���>�(�6�C�x#���W&�k�V�,ޥl �Jc+,'r �U ޒ"Ud�j`��{3�`=Q���\�M:ϟؙ��\L�Y��/hѻ!��-���g]�4`qʨl`��yNH��Y����l�k�-ZY+�$!��O�~�34k��/�$Q��}+M�B����8ŪUG��-0�o7cId�I�65?�G�f��G[9�f�����Y�t�:?��2��R2�h�״�?]���(>����d*ӣ����H�̡���
�����!�ڧ�=Zrm�Y������60�}_rY-y�|V;��ϩ?�O�S~]G�Z��S7�F@=��u��E��r�9�g�߰𡿏q���-�{��XL,��O��W�vl��{1H
�V��U0��I��8�P���T�qN<%O{x�x}T�r�b��U�G"y���{u�*s�iD��*�1;�����hq�BK��$'(�ӶD-|�.�Æu\�����նx�OY?3;m>_�Z{+m�_:�|��w���y�+s���e�"�U}�k~��ǫϯ����\j#9O��]��/Q��n���3QN�Ρ�b�L�ҁ�!���O�<:�/�����	�����:�.�8y��Zfa;cvD�+����y�S�������i�5E���o3����qX3�h�1�r�|߶��2�¶���/��G�[Ѻ�E����<�YQ�˦6����}�(�b��n�dYa=�Z"� �O���o�$.�HȲTݩ���4Α��v��#z�ċ�nM�涳S`��Y��� UM!��c؄�� -�{��=}E����������ɞG��H؈�o��ٓ�����>t�"���b�os^S?dI޵��p����V�)fnP,jMbG�V?�rF��s_���A�y� �؛�FZ%*g��p�nxy��%�O�D�I���6���Ҵ����7��x��C�H&?�-I|�37�à&�d�����,1X��z��(;��0�C[�%%/�d	���0�˶et5�>��ǆ����㼦� ��-?1�R�T�(15�R|���^�����E!�F���
T���3 �{m9A����K�?> nr�;����������ZbK�V�c-�0��g�"�5���ly/S{��#I��H���Ol�� F��v���f�%='}�sK&��{��G�(����txʨ�]�cZ��Z:��T*��Rg�w�%֨��;��ʮ/���J�=ʫb��pG����نr����y����堗��r��=G��.&+O �:J����تc���闏PK��٭!_�Npۦ����^[ա-s0�*�9[ )�ܻz�Kk�"��@�|��EO\����	���%z�.l�)��l��� �A �� {+��&�x`Xe#�����SQ��)�,�i��_:j���>p����LA	���_M�KᢓMk��y�a�	��@����Ĵ�07� �Xdy��az���2&6qL�ţ�B�{���W���4� c�/�˞1��gQ�fb�m�d�RJ��.0v���:���D�annm�韰i~k
��#��$���	�9CS��+{X�';-�t�6��C�������"hVA䧍y�;�TH��MZM��36����p�@,�	,���D�fKx�&�N��.����5�M?z0�Tp��[�X �ǜ<�A�'�$'D�8�˟Y�ȥ1q�I�����Θ����'������{�k�F��!t���o�Sx�	�O��<ߞrF�i��v�S��S'�m�td����z�?�<��!�`C��=�(nS�a~��8n�:k�1e�n X�ܭ!!���	��8~��F6i�Qn�r�X���2�:���]
�U���~D`�`��̵5�`��R2�����<ob٩�e��ع��,&�\5�A�/���:}���K��݅_`����v��W���Or��l�`�4��R� ��*q�݇f$k0�D�� ��J����=�(�|˱|Ë
��.�cu��$<7WWn66��B�f�������5
��q���7�%�0������L59�B��������ޑ>�X"�>�������YN�H����)/�4�OkZ�q=��s��%�.v�<���?�H�����7����.
��-�u�8\e���}K�MM�~��������i/oƾ�2A��O�J�YR�!R����Z���޾�jDgA���:h��T:���X���7ΐ�xH��e	̙��,dc��#��8=nۏʂ駴���;�$�nRT,qxL�V-;j��om>O��{���Š;�$=�l<�0.�8����W�3���Ȑ��*��[�-�n�m��=���L!c�^��%���ʙ+l�(qQ,��,.��2��<�9�?�k�8���r�����ɹ>B��?V'�(VUTP��cE03=n�m-��E��"�N}�[�V�=�pܶ�u_Ͻ�&��r[����/s�ÜA��P���*��c9�~㉰e�6�JEٽ@��De� j?���%�k��G��J~�Q�'v�0��2M��y
\�z���e������lJ�6���_
>�0c�h�&E�`E�S����y3^s=�.���c�~���aՏ���G����b爲��:j�@�޸@O1��hNzbl�:��O�%m��"�����;��mܬ3 r�-)�+����'�5��K��Z�.�?wy�v%~M�B���ʪ�:�t���[%��#O`��ӯT�a�����K#ucaI_-���E�Hy�)��R�|{�W����ԞS�㭤9�s�@��IAp���c1nmv�!w�3I��Z�M�Y�"d���nV�Qݵ((I���Z����������D�P�"��Q������Ql�O�D���)�h���f ���¯ɕ����;{����i�D�	�v�Fk�[�(��ip����:֘c���Ռ!{�P��1�x������fj 22��:+�T�Rj�����k[a������#�Z���t��n�X������8�~ӹ&�i%�����_��9~�r���#��܁$�(��J���+|�eJ���t2����DĻ\�ēS�pC�;'��o߮y���l�jo���F��J�pM�D�,�'�̑GK���;	y9M�<��c�h�(EE3Qj"�uOk^]./*u���	�v�m�߫"O��NR�p�<���qc���p���$����Ֆ���{Oluº��3���a�l�F�,o�4-T4��-��T�"O���ai�5:>#I�����X}��_ �x6��^�9!V0!��Ɔ4{��S�?�ku U��%��v��  �|��2�����EJQo���[��R�`��n��Hh9Ĉ%ն��K�~v�Sd�@M�9����0��=Q �hI���� �$���@k0nhrw�u�P�;m1F|��n؄��Q(!1�ʀ�D�;���'�8�Q�jT'��G)�	eJ��|��Ѵ��w3ے<��]�G�+Lắ �$"> ��	o��z����*�*I*�N�gP#�����*��	�PB�uTC{�$��V���񋽔$��0I 5c�/$4��-�]�1訴'\w&�
�?=d]��Ũ��1��|�&P�h�+��+� ���]�\����I�G��Է�RUW��������(�)sv�¬qI/��jz�^�����A~�Gn���f�N�p�ۇ������85�[�{F����Ć,�'#��i�7b%'��Q��>��v��[Ɣ�n�=i�Y����8�AbxZj�):D��O�Zb�U�X��鏈(���~��=�Iy+�,N"@�5ݙ����xܞyW:��D��
M�kl,0 �Z|U�� 4����)7�w�D���^�'���/_�uxJ�&��� ����Ǽ���N����8F!���R�=9�9�l�_M*��Q.
����HIy�s.���b���P�lg����5�G�?
V�Ŗ�,Kb���&��|��.����R�0��^9`I&�
2����b;�l�T��R��Q���0V|�ks�!��K�6ך4��s�tc���v��6������Z8Eͯ+�H:�V�d�ǋ,W�h+�_�2�a���,�UGU�U���=�bȪg�95�$/b����N�~z�n�����I&}�B�G��t��=̪��L��/,�y�!����?AUx�O�q32zА�����6��c[c�K]U�E�����i��'ǂ1ԋN7�6�>ߐ�߽��#(�An�t#����8O��p�z�����	I��zrx��m�� �Z�ǘ��9|��8����*/qL����Cx����兀�j)��q��U- bS-r��#@��s��¸����$�`|9XB�U�Er�	�����*/�~�J7S��3��"�����ټ*K��� �,�?R�f(E�G�5&��<��}I��p63�@g�*��Z�6���n�
х��9+���Ի��&�����<������k4��R�J�T9�ĸ�\��k����ٝ�P~�"�?��������"���Pd{�;��mD�5� .�����O-��.���e��+�7������U�yL1H�8W_Z8��o@���KտoC��/ 2��W�<��3�rd���D�1�̩(3����p��6B*s v֡�!�Q�.��}<G`N���{���zCd�!lEk���RA���m�r)Q4N�{G���y�I¾YAO�9��W��6
�ҊX�Qf�S%盧�d����2,�i�[��^���|6Ta��\WQ�'ǳ��":����,�鰄���O��f����a�Xs���zOs{B&<����U�^D�S2[s�l��_��{��7!��g��-k�z��^܄�J̃�<�}R<�w�9���>H����$�cT��3�&���tƮ��[z��nT13H��w��� �Ge��Y�8��Z�؊�s�˖���^-V�u{X'��`�	SK�Z6g�b��s,���e�6���<@`OB!�0��=s$�?�dZ��pe(̯L��%pm��g����|�@tx�)�B���f��~�=d���;�Tۮ�#�uYAhD�8��_'�Y�Z$t*m�I�����8�%	-#�IڍOҫ��A�����	r�s�|�)o�&L0�w�'�P'���X.>O�c�p����%S�������	�1H~���\��Y��#=:?�d�"���<��>q1ȋ��2ݾ��81ߋU_@�Q����ww?�j���u��g���:�i�el��6E����tot�m"3�	��S��Lö>��>yH�*r͇BO6}	��]�!��	|� �i��IEF*Z��r�x:
�Ěe�b���-�Y�;�V~W�HC��QG~�}��Ki����	�����8���m����C��t� �E��+w�;���^��P;��$,�]e��;�J���DP_HO���A@������|0t-�FF��S���x{_`'	��=F�Yxv�\������45�$5�ŭq�e��TZ�'rRa\lhk&�3*�i��Ra�S�\��7c�X-��,��y�T,�e��m� ե�%j=9��]���B8�
���'z^.�M���a� ��xJ�4�����r���  ,�d����O�2���JU"��Ġ��B�f�t*�|� ��,h����W�x��mG"jˈ�@���E����nf����u��F���xJ_P���+#�ӏf���{��3Z��w�b3�6��h�ʾw��#jqc�+�Y{�RW�]�a7�>��j�QS��F"0Xb���Rv��K�E"���Aɟ�4o�M4����B�[���ħ��u<��Ul�*��˥��p��֧�"T	z�3�S栩�S�r�Gj2�m���J�h<�Z>��	��)i4�>�tf�����Lu33=*8��\oaVU]4�8�~�9~%���/�vG�j�x����.yK���$��|���hP�u��T��f
(�6�K�[k��C۽j{4}I`�.#�F+��0@��T���_��nY����7i2�t�í�0?D��pvƩ��/�-j�y��\J������,9>�R)cT���m;%�r�V�Y���@I0���E�gB�f�����-�����B{h����#2wE���rL�~�=��� �X��$��D)�{���.�p-s+t�C�M�#�,� 	c-�Dk8�yi��=�?����a����aL��Q����q���`�we����P��������p�l��,VW�.���R�l��ų���ۏ�|ޜ����Pbnn��!��
�O���^5���nG��"���G�k�J��UW�zQ��7t�.
8QF�&��f����p�sz:.φ�L�+��!M��0���	L��?�M*����y��8h���9��>����K�p�?��hO85��@�X:@N�<����E��Bz�FN%K����$��O)p
e�;��zx=i�L�/�w����u!pͤ�&�N!��!'�?,�X�B���hU�_uHj�}�U�_H���╮�!+ J3��?����C>�^P�)�,D��Z��1�"��qE�&q�q�h�V�b��]���聾��h�f �����c.w�	/�)�^��na`�d����-x�F�r$�+�m^�ڹ���|Rz) ��)Bj>t��E�A����^w��l�����
�3�$�c�(we�=&gG6�VE9��G���$�
����;K�Ѳ<��iT
p�>��\������+�"�l{����1�s��~e�qжZž����9go��K�fЩ��������!됀Q�}��tZ���?��hӟ����,Ф4ʌ�a�W���]����x�V�/�E���i����ǔf+��W�Gð���`�Y4T�(]3e�r�*�>0�JV)�[w'�!F�R��L=
S��
y�@/V*d=��g>#*����{V`Q�P$�J�7�V9t�ݯ����0B�ҰӱG����$�E�ƒc?oWD�a*5�-�g��Ϡ�ŗo[@ќI�a������dݍ���L��7���)΋Y���35�V��k�ͭ��ҝ�6�:�0�J�Dp�>���ƼFN#����9͖G�gԬs!_x�]�/�Բ�)�ٙ��,��;L�[d�Hm�?f?w降�|�{���o����@�F�6�����5\�~��15��J��V&W�KS�7kF�8�`��vw8�(Ϯ,��{�Ԝ�������Q�BkGQ�K��D����z`|��w1^ٖЎ�)��@�K��F����@�Ħ��:PEP�)hܜd�	@�$A�<X@/ ��֣�e��^�Ӓ�W���ϢT��e�+б2!H��nlX4���M�gb��1F۫�9͙7-��T��G%:Z$�)�&�d�k��ZW�%)�8�`���R�ܵ��EQF�Hj�z���zϿ9t��kl3�|lo�H��̨Ǻyp������5u�ت���*��7���b$�2�E"������k�tY�Ga�M�t�PNv�q���f _�X�
�%M�X��j����1���!DtMa/�e�0U<�2H�Q]i���tNؓQ�F���2���-(z�u^E�,���܀�''���}���_h%P�����d�2��Ws���0,�*�T��e�i�Rvw>~���� D��� �c��/��4*B�հ#��IO�ׇ҃�G`���T�Q��sƦ��d8f3�ɐjH�Ca��ǥ��������t4�}|MC3Nt0�#9�̔dl�����SU,С���3ibJߟ�JU�2�/�\��A�l'9��]K��-���d����]��?�os�4_r������r�A����,�t� �C�kj����0c��rNow�υ~x.��ُe�<���Tuu/YE��i��_��	�>/*")Dy�^����:,hEͭR��
��;�j����B��i��Ѫ�<Gp��,҃ �^^"?�ՎD��+��گ1����n��=�>5��4��@����`4��(���9����'���`E��k{�� ��R�!g�ð�@=���5pd���7�JZ�M���#:�W+ �UQ=�k6;�k<�q4�n��!��mޏ�9���G`�S����2<O�&R�c�]�G$�t6�.r����\���@z��43Í��`b�:������.YE�����/~(�SM��$v^A�������Z'^��{�c<��c���F yF�@@�����nԭp�������o���(M����Q�$��J���:^v�/Xe����I8H�z��R6����_W�,�"َ�P(���9��L���e���G�jA��|ĩ�C=�3���\�bp�'W�4�l�&��E�oI	�X
;�e,�C_�{�������u�rs"xô{����(�v���Ôk������@z�:�,�Q��K<R ʸ��>��S��������*ְ��ͅ,��`G7�p�Q����@�t�Z�_`���C+�W!��
���7�����x���J�V�D�w9A�u8X�*�m��!���e=�&6���ɐ�o߆:�2��ɡe�J ��u�&�Rw�e�j��J0�l��P�&������~a�_3R�e��X��瑎]�H�C�uLφ_.��h�ݎ������D�n+��K�w��)%�wG08�vC���)�H2"P}<�HD_���,ff`Gz�򲻜�������ޗ+_�l�N�aڶ�.P]aa��M����Įl�,\����UY��'o��0% ���q���<R�$`�j<���a�쵩+H4����7�������}w�VE����v�v�[4
>ёtZ�"�����/CY�ٺP��ZY����y�T�ҋ�=U��Nڴ��o\:YF�i�EW$����-�.�O�"�T��JL��Nu�F��L��]x@rR�Eg@2�
���5�����}�!::r�E�]-GM�`�X~�T�Ztఘ� p�\� ���.�5H��4�G`��A�"�rDS�?���aP>��Mׅ�N��6Z���$��R~2F ǃJ��d�a��|3�*�nЌ�P�p
t�&�5t�td�w'�X�0A�E�|�jp�I*��]���۠���R.!��n���D���>4
�ʔ�M�'-yU��"<Q��t��mT�����,�u�j�%�֦�N��"��y�<���l!mh_&��0A��v�ҟ� ũ�;����eu��h#�_��ƀ��X����d�<�"^R��bV8V:t���PP�;���[��Z!�T7GD�c &�F�3.q,���C�VgۂD�q��\��Z�"���PE�Υ�O%y���7�}$&$�(�E�=L�߾"���F	a�G@�Eb_\��fI��J��h���w�)�6Ɵ�;�92s}��\C�/�j�?�x�I�p0�P��!�|�.�{��Z/[��0ږG$���F�cw.�E4O8���z�E�:w�&�HlL�M�60W������Ҁ6, ��%s�鋀�Ơ��YuIO�}d���n���E�U�[���-������۟7��c�(�"����b�A���od3������*&�q�t�_?�G^\��&��f�˖z�ʝ~vV!�5A�-kb���K�6a�=x�����d�0�GJ7\5�R��qTh-�HKk���4mx5<�5�T��i��	�<�d�]��F+��с����׆���#���E���̹��h�.(���FhRn���5�3#��e�v�MA��lK͠o��j֦��[���'�����5ZṔ E�<�s��Gzw��{#w//�P�Lb(?X��W�Wi3Z�x��~�.8ɛ�S`��l�K�{�OXi�[s��� �Z�N�~D�"��7���Q�m�Ҵk�X(IW�dLej�h>eR����R/����}����`b
�|e���G�c אNlѤlD�cA%����x��ãtU|y�5%�q)PY ���<��k�v�$����;��R	�xc�B5{�BDJAn��d�ַn��;>���|%����,C)F���"�U����4ǫ��O��r��z�a���U������o�$��e¥��2.i..dk� n���Ο�ԋ��;�����kټ�r-�l��"�W�=�fh�M3��9~Uk8lp("�zC7e�v��W��\Jf���I8p�(/e�!��9��d@W|3$BLj��a��Ѱ�����24A�C�������J*�,b�}���}�I�zAj'�{v����B5.N��E��~��tm~�4�[�{OC���)�$#�̘̘I&��8W=/�a�75d��
��9���󐷽盳**��G����ip�Agk��Z*:-oJ�EL
�Q��cR�&grc�� r=�2���>�*ݪ��A �ȗ�-��{��c]�o�'���\�e�j�I)��(��8gdCV�sq��n��`3�tb���>�d�j�Y���=i��~���N��B�-��.:�����fx�Hd�?�8<d����f�C�8�0 ����^�!�L>�G��?I��������c���^ۅd��	$TJX�g�]

��)%�����B����b��E�I1=�S'ޤ�{`:�6�5
aq�H���(�zy��������|��iC�mu�\z������3c��x�E�1�Q���YY��\�5L-�>�f�Y��)��������I�C͜p�K:cR̝R��d��%�ՙXqȩLՎ	���	�B�pA�� �+�ê9�Ti3��;�#��7�y<e�0�kLd�d�#_4���$�cv�����E��.���՛� ��y/�F�m.�҂��Bwv�S���H�]�W�+��'���0��L�d��v���sϥ����ͯ2� ���d�Ʊtdȷ�lxl���d��S�ED-#�աC_.n�G�����.~����3Y��� rY��,JU��� l�5ƕr�C�1�,�ꁐ��G�����1,?�]>�|�iލ-	$������o�\$�7rC����x��`���	h	�� �W��ڛ�T�{/�Wh�Y��2���\�&�3���,�+�{a��ȝ�n_���Io��R��Eїh���61����7��JGd�Ha�������ڿ)��i1h�H<�@5�g̹�P�>��㬍b`w�O�/���2�䞴@2���p2c��Y�E��"�����R-ᡛ��o��D���a��9g��Ĕd��Nb��l�u��'�a5*�$�~b4�J��G,!�f�;�hWT�\u=-*ݐG1�'�H8���X�Z�k�jF��������o�ڽ�3T,����-l�'��%ME"�g�֗U��v�Mns���ah~������@��Mԕ�"�F1Z�_(޴iU|9E��To�	I�\�9`�pc��H��<Ç�BbO�^��G�a{v]�*�ռ���`�5�/��M�2X:����Co�c�w�&����"-&�Ҁ�R�}�U�T��aT�XD����-�#���	�u����ƍ<M���B΁������<9)���ҙ�Ǖ7V	��l�8I��"p6�Q�TPtOԜQ��g~c����>8�NZ2#�B�@�^�Ƴ̉�q!*����K���0%+��U�B���ɮ|ɉ�s�����k�T�7����e+���M���!Ë�^�4XUX����Ψ�PRPBP�(`}$�7�δ[��Nom@���:�LW
u��bMu�i��$It	%̓��������5���\���������:���bo�	Ȝ*n�"����co;�g��Oo�O�]cć\��g��st�!�k'`�8�P����!���������|P�}���,����6�z�<V�U��Z��9���Cל��`��6��Mq�.ՁLg~0�FoJ�6���:�@��=�'����L�$��!�S&��@ٷ��P�9��>�<mn�|V�&?���}������Y��A���~�L/�v�J��ݔ}�/SM�X�[�����ad^VI��<���b�����O�~�{�m�|6�U�P�m�m�qi��!lb��2��r�Cc~y�A�`0t��Ar��}JF��7,�Ă�.J�dcֿK��T��͖#/�c�i�`��k���ɤ �
ċ�j��DZ�� 	�[��5��CrA�<.�=�n�b�@R��P�,ɝwI�zK}̖���جP�!���[�s8�{�[��_�����xBר����GW�H�x[~�^Z���>/���l [[H��~�.�6�� ���`�+T �V���6Q�:ٕH��d�������*8@�Mt@\���q�6l�� i'���:�����,4�6r��;E���#�uƝNV�D��c*3���hڥ���4e�['u���Wv}�6�-@~�~�{Q��s�ڱ�+�z���t����:</-���:����D,��<��MZ� �A�
o����?mY��W�l���	�Ue�k=:�(�a�9��ZM���W�ђ-[񐰘?���Æ�����F�j��Y�b�|1��O�?=4C��F��.�8H���7^~xXQ<�e����#����ɟ�F�jX�t�K�υ��JL[ti
�5@�q�
��J֏�,	�����.v��R4C<(�`,$�ρ��@���iK�y
ee
e�Ml��`����z�K.i��3��;�	ܵ�A\ȡ[�=2 gHw<������M K,���1�x��i|u�.�`=��l��C��#�3�>�b�h1����GP0̑�Fi��U`�ج��^�8���M�fS��.�s��B�Q��O���{$=I�nt��PM��;#�%��O�튝�|S�I���w���_ū�t*�77;o���A��5ɢFGw9��E�q��@�n����@���u��7[��t<��R� >J���P٧18}sV�
N���I�6��OI����L�gU�v,)�v��7%�l��|�0���R�=l�׉���#_/R<�^�/qXp'���)�0,qDX�"�G�UӬ�P����Z�^���nt=��=�b��l�8�]��U�
�U����$ttԏHV������/�\*�*�&�(�F���u־�)�Ʋ�wɅ�Y�2�������-�OvH�����I9����������٩�3R��8�O5ـQ��ExM����A�;�qs��3]H�1ǵl���'cu��(s�VѯX0*�+��k(��f�V*��!����gR~��'�����NS�`P�6A0��?	[��|�?��0sO��q�{�:7��;Ud21��i
	S}9}���UqU��@r�=�e�B`h7��7̅o�" .,PBౚFu�v{����;R\�<OLH]��J�F������N�v�fӿgs����|͇���V,k�^F�s����GMD2]�S���
m����}��W���$�}g��<�G��ѩ��[$FW� "��hB��G1��p5u_�d��c/�� ys3��g�ZM��0�3��+i �q���9 �)+�&�˛��Ѣ�U1�L�b��o=�O�d�E��GVD��u]�X���{��b(ש�>��d!��u��d�Vg��I2:vU��^�~Q�T"�)��h�~؛�A�Z�^L/j���r��u�c��h���3�o��S�ؤ�)`�b�Q5_"�ީ�<���G��\NDt)�s�����ߡw�@I���b���YGp�q��*���5����ͥd��5s�ذ�zkyV��z�.z-+�� U����rU9tlnu~��Z������;Y�z�3qӾx�=�(E��"zE_JV�5;Y��n<���d�S�շ���6�C�R�͹���z�np�����LV�ac+�^�A֊���/\p�*�}f���	^-�C�(9�Cd�ܹ�6�B��`�Tat���^ȏԽ?5���m�e��YH��#�c��p���ͭ � q��4l���t����>���#��p'w����'L	Xh���lo�J���ijs��i�ߘ�"W�C�wXoz�v�?����JlV	�Y:7W�B��e��� G#0��b�}��E|i/�	>�4�Xr
�s�B-��t0X�I)M7qYVp�kAU$I�?-�|Ѷܶ�dANt����jS'�y
[��^��Ɵ�jmѯ��=� L/��ʟbާ}E�Jv�8�����r���~Vc�G��Ɓ
k��f\��O��W�X���p�n��o<�$�l]�abkŚ2r��.X_��j��.T	�H�.������Nb�vnyp1b���)���.އ�=}e;5_�d��;G��9UCTj���p����}5`on�{S��� Lpڏ�@��,�i#��V��Jo�ZJ6��x��	����p:,��8��3�B"���}c���H��7/|�8��T7�7�g�=�}�#�oO�c><�!I�ó�����S�U������+|�@D��8�-t^��-�"�[;j8��A6����+5���뎈�!��[�Vl�6�P��rp	�s�,��u���Z������B,wϤ�ay5�
��6��!�e`��v��	��o�F?��
� D�'�P�JP���`�E̥?�h�(s-���,g�O�ҁ!��a=�,!B)��#H{��T�~ngW�,[Z��U��iM���!-�'�XYV��`a*?7����䀳�S0��)j�xƣ��*�I��������A#"�M�[�������|��\9m� B�҆V^/|�h��[Ԣ�ÊA��ۛ�"�8�<zѕU��L#�%�o�F�{^<7�e�x�CԿ�&d���W^�\4\��i�N-]T;��Zp ܠ����uMj��j���*xLU�T�h8�1-�p��]�Z�j�Ȥl|M1��{e�o��M�
hhݦ��m����[L���F�}p�~��!�֊f��b��o� ���d�2#����wؽ�脃GX{�F�OXz�C�#�UB
2۳�
W�U�=%g�u�2����P� D�̩��5�=�����<���E�WG�����aU0�d�f�����^ ҝ��#��n1i�O~*ۭ5Გ�!麈��$㥼i}��XvCe���
C�ˇ�6-F�$���w�m�Y_���ciI���>.DљZx��qn��/+&���\��T��Mj����ѯɒ>�l��~�AT�V�F	�؍��B_{-��ܵ� ����B[F� ����Ĭ��վB!�/]a�P�:��r�ݖ��sTc1������8�,\hs_�{��إp�Ȑ��b��" ��9D]s	���n���o��ʲ��w���0[��fc��zS����R��3��,��iy#L%���C:�Ϩv���x�����^?�תX.�=̷3P�s��}�K�$���%C�f`�)��l&�!E8�N
f^�7���1՟c��2E#���8Z\��+�?<���r�#�@�;�1���U��M�D܃������U;�m�7jI�qB�G�!2�|v�'�d�,O�F��L�m�
�����R[��2`G�Q.�smIfba�ĝJ��ԓQ	`5oH�3<Q)�6OB��D�q�-�Ah(_�
ʼ�#C�e�`�+����ܞ�Q-��{�&�_�\�b�팂Jc[�?XH5�>�'���(4�z�������>D�+�f~;����Ԃ���N%&eB瘻�d�ԟS���;�t������:�s}wqi�n�n��z:���/,���z:��@��-�`r��� ӧ6�z?��-��j}=�n.�(.��"g3%h�i]���f����N�U��։(��Z:�����ֿW��y���&	�P@�Lad�����R�n�A�n�I�����5���ۉY�j��O���A�HT������a�c/ph1�C�	���qmg��)����ր��*�����<6���فG�^��r��c�J��/����t���W��d��� �؇j��\��i9� �w���5��+�g֍�pr̨�������\�od��QU�>�D��l��ٮ�3-q7�=d�^��4��Z�o�ʘ[?�h�m�)�k�S$��1M�c���<EF�쐽],n
�������gۅ٘���؞�WpyL�������\D���{7�����@k��\S7�p�r��k�`?.2�1��4�m�	��A�ڈ������
���\����a?�3���&P���+N�N�bV��^�LZ����#��;ص�Ɏ���֟A�w���ypd�sa˃��ڽC��s&���֘�}Y��=*�5|�X��i��ש���z<��B,�3���	�>���I���X*d��F�y~V���ޗGb��0_��D�5�F*�!~����ㅆxϛ�M6f� G���p�g߶��z]������*%NRqF$1�|ᚷ����Fg�>��L�,��@"��>%V�f��$u�a���=p���c:��Y�@�Z���e��O3�o$c�T<����e����{5۶��륫-}��W�ݓA!��ZR�S��P�l'փ6P���g[�svq�~sC��/0�Aů����AC|&��Y��dKK_�������k�S�����k{:>�_F�T�������Dw�K�YZ�`����k���Np��k8��R�`���j�5#ɬoJ���{�Ơo�\�.aa�'�v�؊ߗ=v�T@őe�i����pe����p����RA9�y/��g��R`��`<X���A��.̓~��4Ж\�h�?4�1-Fbޱp$ ?�y^W�s����50�8�8R��l��׈V��C��+��c���I)k˖9��.�Mԓ���FXFc��{�}��G�M4M�|qg"�n�#�@�%$`tc��U�	N�N�k[��(�֏��ۜ�X���s@x����<���Mh�4b�"�n����/�E ��O6@��"e�j��;i���b�w5U�Hi�@B�A;��y�1Y��Ha��K�5�D�E�=�#���>�y�pD��9 ���̣ƽ��΢9r5j������n��mH�V;GpV�q�$�|8��
���F�[ǡ��Jy%9^eɈa��W.�������d��I(|J_�`}��.ia�kX���,+
�#6�vd�R#��KJO!��@�M�g�-g��Y��&L�T��D3�z\3�ٗ�s��"������t?�v ܉�H�ULS�D�3%q����֥l��<��ëU_$d�c��$%���P��D_u��[y7rXl���뾗%�&h�?+��\6O��n�9 ~Z�tA ����Y���5H�;�M�!�]R>a{9L�<�O�Qj+�gF�fXa���ݔ�����l��R82��?#�Ax:g����C�#���%KU*S�g�v����0�VS.o�sW!i�+��W6���R��u���A��И�C�����5����@�����:�c(~	R.j�,	�B-XTB�Ǖ�4�o��L�u��l�g�-�=�`Y1}��<�s�ԙ���}Ľ��d��_$���hz���sɏ�<4�Һؽ<�+���^�Dt;�V̬8�|^�V����h�����
b'�C����r��I��#�TeBt�lI\8Á�)$�Ԥ�q|^X
�IFw:#õ٧W��p�	�ɯF�z|��l�K7R��/��s��PqF��Yh�!�>I��nUI�E&�dG!�k"�Vd��$��+�}7�r�4[���؂ bޯ��Y�8��{�v�pE�04H��O����.��cE���G��A��mPB@wG�Q3yz�O*|A��`�`j�T��1�Bk�/�_�6�@,h!f=�p��A��NW��3��*m�s�‥H\f<�J�w�:��M�CG�l��������S$$�c`�[˗��d}؍-uD��J"������
���mZ�bkЕ�ڼY�[��IԐ�fy���p�6���3���Pp�.�0�ߞ}��N�U�U�K�Og���m�%�6Bq�t�~<2 ��%�㷵�>��Ɵ�Ja/��p�^��2_��IME6�a{��-&��p���[CA0��_�F��m2m=��z%�.'� �\_��E�W���&����\��I�����x��6�Y��^��D�� �*���ps��d��G-,/��6�j�e�� ZoVq�k����]����YI��)��7�`&ӏ}�l1Ì�p����������p�폌*����ր��O�ØK��Qu�a&�@���B��36��]I�ty���a���f"7M�De���`��$&ń;�TZ�j'��$�������\�B�YՂ���V�ڒ�"��ϱ��O�����_�IgIC��&*2x
'a�}eKl�>�<{���~�������䮛_ނ=N����L�$!��?�ﴹ�3u�����x��hg�4A�?M5PY�֑M��oqK����'���@ľ��h�n��%7 B[BS)D[	�l¯�N�m;$�x�_������:�d^ɫH�W����ä�K�aZ�Qʼ}��7U�K�E��$p��ewb����� ,�U�x����V&)�(PN�f�r=��`?������
�:���? F�?��-p����d�hv �<<�y��\���##���]%��>��`��=b��(elRf�n!4��Y���ż7�nV��C�;a�T���r�Ν:��)�3��Q~%�t�RZU$t�!Nr6�Im�uf����Ů��t*ry���)�wBɞj��n ���a�XѼ1�����v'(���gD/�U�	L�������w��_Un���0�7���_���������4Tj�M9���9�-wU=(s�ڲn#�e?O<�r�9\k�s��_I���b�+슾�kof:��!���7�;�f8���.�A
q#��.�#%yb'�0����|b�:�������D�S�C��.��o��ܭ��X����P|��ұp"*lmx�̏�Q��<�p�q�(1�Q4^��.w�.��1�H,r� ��8�,o+���x���x�,�fƖ�d6��na89��6o��IZJ�t�x��h?G7����'נ���-G�O���k�������h�j������� ��2Jma���XG��Dn&���e�dnI�I'�@�X�%18EN�i�~'��T����بj-��g(+�[�:}ձ�����%���3�oo:##�Bt<\�%��/Q�[��v��ޞ���Bܶ�qE�gK���&0A�����o��Q���h.�l�Ri"ȄW ������0S��	�Z7�Ś&OkԢ$��3���|`����k-< w�3�T}�|q]$b���cV�Ќb�������ą_�tA��j&sI����e�����3��=�w �`9ϰ����l�@����R���|���U����3������ �
�<�7���9F4y���3`P������	�!.z<���`���y�}NVڨ^�ޢ/�m�n39'Vg��iOב�fJz�p2{P!�Z&MA��+W&P�Kѿd�Q�ެa�c�b�������|yj �>-K]����f�	j�{� ��2�'�Ն�U�}�G"�0�/̜���M��A��Q��"�Ը��1���U����x��ts��ඌ
-��Q5�	��z鮺F;I|��
��U�/z!HU��x�QV۾��U*I�l;�¦��O�d1فcg�ȰϗYU�_�pq
�����H��,�J_r�ݬ�sc��R�������l;�����sW'�+Ax�Y�]�a]]"6�����w�$P�b1Xrg����������*�׆���쎙.}\�����G�JS�<~*��P���e\�Qަ�^�nZ����N�PW%����ª���;=zh-���'/�c$��{�����xThİ,�d�wt���*�e�.�u�x���%��3�����m0v��� ~��$���O�͈+��8bF@Ê�09���>Za� ϕ�^��k�!�ΰ�y��Q>��M��S���X�T{v��{�7����pn����Zq�C����_왨�]�)�IA,}�V�
�j'5���z(VI:�z�1��e~��L����q�
�Ag�v��$��t��m�V}w���i1]�G�i,�����|[/dw2R9b������e���8�a*0L��C�'��L������c�'f@�z8�ֲS���Ւ�7;�.X�A%���)�=�ٔ>~QJ�폹�ݭJ2����Uߝ�N�y�`����P�e"�Qn2���kc T���b3�R-���:[8�E;�ˡ�Y
�C�o��Y#ҀS�&ǎq=�g���	
RGFY��!��7e}��߲�w҇#�V���]�c��CƬh�f�����ً�̔��f^�+6�:�"���
 uv��ؒ�y��"6Pߗ��6�n2e�X͂!��n�T�I�$��Q�d��	����Dq7h�!F�4N��AN]�r���Yצ>`���|�p�z_� �_�2V��Cf��\8:C0�������6��o�����1Z�h)�Ƶ��5g�R��r���k~�����n�M���Pc���u�w�"�9���(�6��V~l�[��[�*<]F���iys�7�
�()���r���
vReRV�t���
(�l�D�T�Ν��bõIo�C��ú�m�� ��q���P
E����?dM�ߣ<�Ld��G1���B1Gi�%A�q�KB�����㛰��"d��2N�S����.x�
�9g����e)����H�7���"2��ꆱ��\ݳ�ls�7���~߾�z>�=4{���wK��h���+����Vһ<SGP}�$U����� �������lf��6�Dfe�"�Rw�7����|,7��
3x�߫=�ي���/�U�ٙ�ؤ��6��QG�4<�p�RY��T����l=�7�8�n'UlDp+e;>#���y�Q�m��	�����t�Y���Ħb�kd�B�����������b耔�ىgM �l�~SO�Du�5��ݞ8-���~��up�?�L�:�%�r)�w��i �_�[��>�S���U���E�c��;@��.�,�[j��a.��7U󼔍�϶�\�7�\���E�\lg���]�A�[,�2o<�Bx�͵$��݊��w��	����ޥ&E����wb�cp�
St��N��[�����踓QB@`P�H!<z���v�����R�w3�-��>)t�m�$tꗼY�um2 n�*�&�4� �_���.OX�T�ѱ� ����J�/�7��}l��O�Cl���Cڕ4.��)u/"�3�L�h���0ڹ:5<���i�9@�����H��~7��_���g������5��{�olv�-���#2E,O�����މ�ZY!�x��4Z1�kBc]����!�,}��$��aZ$��G�u��|�����}�g#���+R�\gH3(���,41��!�}h[��᯼\��C�����OB��{�$:��0���Qs3�;m��ڜj8��� qTq�蜍�d"4�z���1�����)t�9@	W�5�|���8���2�Cv����C�Wt�X�3�]C�m�o��.�8��?����lIx��
�a���T�l�il1vR��:0Abh`��\��W��u���P��лV���$����S��4��ہ����E�$T�Ik���tW��B7#$��]�[p���59�F�'I#~�ɂ�e�PD�xh�5/��C$
TA��8�>&Wq5R&�LD8�'����ŨυC`�$�X|&ߓr�k���@q�����]�i��8>���k|���r�i_�ֹm\��nxSArn�T<��&HBbr�Q�fa�¤	�"�R�ާkn[41�%�~���Ќ8�I����C� @SP�g��~�$))�]����C��\&G��2'��\���rJ�C����l?��P�V�*�ڙ�_�z>���SRX��$�L�M�3�~����d0���ҷ�ֿ[�^=�7%�ѫ��y+#@�͖���7�K@�%�|)��|��~�h�+#�z{Qw�0z���詁{~�9�L9��`�M�{�%VU�K�닲ѯp���ofV�t�B ��K�l����wӪo�ӱ�+[J�n:�8��V��8��S�[�;��#L�>=lS�yNc;�QO�Z,�O��V�;����w���f
�w�UQ��{��⮚\�7�ή*�G�ūi��#rF�m�|�k�ec*�}GZ���&Ό��h#=Ú���b�y��Z�E�֭_��_�յk�v}a{DM��!���G؟�J��A�G�4�^�&	��T.�F�Pl�����z����;��Y�+4RK�zjP;ug���]�/(����b��g�%�[�CU�����C�]t�x�(���켪��l��j���X�-*�B�g��������ʰ�a�� ����o��2��F~}7��w��h��L��v�-O`>�`xFSr�8�	�=\Ŷh�S%<&�H�ʠ���<���j����Z0H����";��[`_�I�S��:���)i���'����(qd�� ���}��f�M�:�O�ó�:�-�1��v�
K�K��+�Q[��O�wH�LE[������Ԝ���~+a�e���t�7H!���z{�8�O���v"7�~��mk��1�T|Mb�7���4�8�Hʷ��-�o�P��$��!��O@5��� �Ƕ�<�B���Y?@���`c�_���K0�]Ax����y���nˍ�З*�\c�T��h���3�1C��@\M;��?,Z	 Y��&���A����J��mz�)Dmo�+N�ҍ�đZ�21�J��N�����G7��S���,����Y����F��z�J*'\LZ� �:}�?�ffw5T�d C(�u��B��5�uOYg�PA٫Z���g�xR^��a����(��v��d�E����i�iZO�+��Y��A�D�Ц���Wl��ֻ-iqiqL�c����l�ϩ/%-)�B<Z����U`��Xf&��mJ��Aڣ�NI_�U�]D2Y#�k\;r�簳vu!t�W���֦�?]zB��yg��Ƴ{9�E�=љ��N<ڨ���'�F^���9�ǻ�̗c�7"�����t�q/Mj�����j`�Ư��wX,�XQ���|c�ً썊@���ܠػ��'�K,� ����O�C-�㌗ߑ0��{Xs�@��h*d����"�C,��c1�z�}y����E����v:��p6F`{�]	��QX�1/!����* Tݚ(�����i��
�.f~%s,���m���?-P�6F���g�/�@����]��"l� j��L����w���	� �ڻ�\
NK����{�
8���%�l�1��lӤӧ�%��7���&H�A��N�����n+Z���
o��)s��|�f!ru��~����l����_����j+�8���0����i��[�N��_��2�	����-�f!W�&3�<�l�����\��]<sǻ�)r1%xۯ�_T�w2u���dk���l8#4���ׯr�LFh�}��A]T��"�|k��M%=��i�f6�R�&d�-�΀��a��&��+C���0��uuap;J ��cw�]G��2��M�/�'\���"�7=�x���I&�����ġ�.�1���VBdι�����Ss����h�l r����9�1٠ �[;L��'�>�����O���W��Ýo�x̵��7-�����6����<�+E#��v��m_�B�S��ZW�X�/�l|$'$߳��sV��_m�6�TƬ	�
�C��[tn���L��;%*���UhgnpʙJ��t�2�&��P�{�p�S�G����4�f��RiXQu�q�����Z��������~5��[��':��'B �hr��
%xT��j*��$^[*꧋��}����v4Rܣ�&����V����x���Y�����$��!$�L���7���:����ǅ�ĭ!�.z�KEeR8�I4�x��f�pƿ�-���h�&�n[�[Ȳ��;a�� t�MPD�ҶLn]0Ee�.V.�������Չ��0�3�dF��-([�#�����r��ImRP/����-�~0I�<�i��r�Y�%#c��Ҹ<mhp�kh���qq.��G}�L'H��Z�z(��)k��tv�!ɕ��zԨ�Q��b�?�myp��������p� ���$���:t���VJ���A����.BshD%��.� �y9�mB7����Iƙ������yh�Zn���e�8Mb�V���f�$zEy���ո,�%ڊ���l6�x�u3}j��i$�Pq_T�9����ꉠ�:Qy�rf��S�o�*?����xH��WYay5���z-q_n�]��)�"9�H:U e�l
M�zm�\W�%3xu<6>��"f���o�����xGR���0���J��)�M5�Z�$̂��5���G;�d��닄@��JǮ�����ݒ�v�������qK	�b=�^��J������u6�#
o��G��� \|���H�����[��t��E��ܯf���}c��!�R㲄s�>f��x�M7�)���L�ܮե��?�<**��;!����r����.�O��1p#�b~ip	�X�u�!(A$��3�����ƄCY�s�*	 -zǋ)��M�G���2'A�6�t |�����R����X��^0��x=�	�A�����~�z�������ʿ�5�5~kvk����]��~�l���(=0 z��)�.�D���/�Ò�p�����G����\t	���m�2A?	�����ŭ�B�YX��Q��_�K����^\b>2�gx���Ԣ�6{R5����z��GT2-�����K�����L�BE�������[�����؂	��h�ky�<�F�!��Jҫx�Щ�t��r����n1�W�yvZc�������*F��>J�i�$����r��T�CxWw�d=ae1��b)��<<`��pV�-<���s�u�&�R2:�4���T\��C��"��ț����N�v`���f�R�SZ�'f`�yf�%^;#r��`�C���yΫݕ}/T�$Y��$+��z:k��>(�_���A@�3�c�֚�)+�y��q[����$!��UTl�ő���D4��6>S{E�n�Y����ˏ��D��/�%Ψ�ҍ��L��y��ח�#���bq����b��փ?�����R��#c�	�8��E�Cwj��W����GZZY�4�z��j�$��_~�;�M��]6B�,�?�L�ϩi����ک��n��B�Dc�l��Pz�#X���t�e��\#����䉈���l�-�veeW7���ެ�[��:�mP�x8!W�<�y��?�3ϷKt����Q7����R��^J�7�� iw�o�����@��Ґ'��}��M=k�C�9�u���+v��Fuͅw=j��2�n.���qe"��W�L��o�ə<q����w�+5@m�ta�E���� �	�p��)�
� ��3��X��/�0��elkS�;):f�L]c��/�d��>;P��R�a�Ź�p,0Oܛ/�w�xOiG�)C�;�9��y���5Ne�9m���M逞e9*U���p6�`�|(A c驕g����'���K�嶔�JU�	�՜4��O7�Y�:����]�@3�k3i�|��v8�rSRr��v�}!�ԃhz���v60R374��FrјD�x	�y��,�^�qYC�nK�3�\.�ny��9���):�&����қb��1[����~ˬ��H�j�\[I�2۽�#<�����Q:e�dU��Yu=&��}��;ŷ�& �|	?���ʔ@5'&�nU�z�<n)o���L�?x�R?�����,.���Ԕg%��(q�?�
g�m$rU`�*%nqh�pr�*CM�[�`����0W���������;Rfެ�U���ߓ���-�����Ĵ�=�ۥ�Ч@�I׭?�*�IJ'�
.��f)^�l��k$^@�tJiB�3;:fBi)��,��H�N� ���.>�à�sa�����RHi�)�>���Xʖi�{ngl��K���>�R	�	��������[��&w��&N�-m��ğk��y�S�@�Ya�rq���+�gÊ��26)���������J�'�X��3C�<O�q�4{1�>����+�^���˕�[��xu�^��w�Wa�"������p��q��#���7�!p�S�彨��F�D�K�OIx�0��_gn���Ԕs<��C":�b�d��J;B�c�6��[X�
���$��%� �\/(o8���3&�9~�D�@����U�`�F�I���$C	��m�Z��<�E������h��Y�V���e���d� ��֘�����ayr�W�\����ˮ_F�j5;��OR(� ��IC��?b��|���$�����`��,�L<�
��
�������;�2kͨB�k@ة���hs��.*�N�&"0P�%ב�b���M��o찡�N�S�K@Л��ښ�ܱ�cY~����dz���	�I���I@C�F��i�WeX~���o�?0ل�P踑�ӴR�Ҁ���?k��m���4IE���ʈx0T&�1�y��(��|Q[X+,�C��x����=攮s��E�dׇ�Y\�cA_?��Bm8��*����!w@U@zXG�Cd�c[L�VF�|]x����y�6�>'�ʀ���s����f��������;X�-=o@1��h����t|�Gn1c��!��B�c9@m�[Dn��>�>)n��b�z��h�5��]`�<�$��^.�4V	l���ɛ�r�����	�4n���P�G�7��/B�[T����|���a�db>�ȩ������>$�ܙ2�t,s��K�ŋ���e-���,�f��$��[��e�.�r�	g2��o�浺"�[5�-��(Cǧ��9����o�IHd�T�УR����,ȣ���� G����^np3 �H���&��:P�2��a�6��U���b}���V��mv��cf|���}ڡ�J*"eF�p�F���YB�	��uH�g`'p�D���B6�y�=���J�T�ɒu�*�Ԡ�)y%pqv�	U��_��"�+m��bx�?�Ji���f%;%�o�����x��~{Z����ƒ����PA׺&׭&(��|�}�z���=���h�/I�)���*\ub���A�K���2n(�g���>��0�U��5uե�.b(�C4��%Y�9�d��2�@\}�ߖs����<��\�L��k��h��>^�,n3�+HAً��z���t[چ������`=uA����q�ت�8y����Ĝ<?w��V��?R�N�2���,8��w׬��O#��c�KVc�xe��i=�.Q
�\5��3�h����35�� ��$�s���oN�bp�?�C�T����;�*F0�"B�Q�N%�0�g�r�=��{{�P���<��������Ť6�kLǲ(<J�kn�oxIZ�j��n�+��SL�?��D�0� uv?�l谋NO�F��4g�#�F�r0��1M=D�O�8ԑ�1Tq�L��;���+��i&���}�<cYϭ�:�6Dxcb���E��f�7�?�yŚ4n�/�D�%�����<�H!�?Adڣ�5?�Irۻ��)a�rx6��r���������S��r�j�e���dWR���7y�g�Ĭ����Λ������U��'�6Uay�8#K@b>�#1�tN�W#[����~	�K\����?�F��E���AN ii�ؑ�ȱQ����,�Ω,n��%V^T�y5�3��&�Aĕ�&Sl�ޱrR��,�R�.�L���t�X;(��`���h'�pc���p��&��\MeqX�ɚ�� EMSw7 �0M8 �p[�#��H��w��d�!����%��Q�+�.�5J��Ds��m%�fT���3���T�|9��wᰯ�V�XЄ.\dtS(ӿ�;�L��1r�:�!��!�ݘ�A�v�AA�wy���0�xm�lQ�]�>ro
��+�Y�]����%��#2��4��~��Z-1>_Z�RW)[J���`��H�t�68�����SG�)��}�t�<)љR:3��Wx(�H|�n�Ͱyh>�{����cM�\�xɔ���klXw��$ǿ���= 5��`�1_0jש��P��?�{nT���#A|���Z�mZ���^�eV?w�2>��f��*�6��)��
+�[E���D�Kt�4�<�=��Y�� �T�;�iPBj`���!�ƿ�@^���|�D�'b ��x��,���K�>�n3�� ZԎ�c�3v�t����g�>цA��l�����b�<�}DYے�!jC��и�l��(�.�k��(Ը���� ���"����;�\K'fO�ӎcS�, ,�V(��
;zE���Y�������|0ĥ�?��X[�d~D	p%���;�����Le��BD���ZC�[�ȈP�'ꠇ�fnF��Hſbu�N$i��o��#r�^�sE�Yfrr!Q
���/�s9��vD����"���y��AH�%��p(O��0�l���{,�Ej�p�"�����YM��O�@�@u	���a��%n*5�^�}��A��Z���О��쭌.(�_h۱� �;��-�{�hk�Y3�Y^�0Q��l� ����8+��RhU˙���_�Ն���6�EԹi_��a/j�����g���#����|��:�/���"�����s�m��ePK3��6Z}��@B�\	���˜��������ZGi�qO³>��䓉��٨E����$���x6��ҟ'��JR�&B�Kd)	:��H�o�"mڱ֦�M!���hԂ<h\m'ٕ7��(�hL��-�g��GT��yڇ.s��C!�D	+5/�1���w��Þ���N���TUQ��v��B%q
dڑ&�m�ɂ�=Jq��Xð-�/K=@
�)�IK����c����y�WQ��6��#T�,9�ߗ�!�ӣ;Bd�I=��1Zp�}W��ߜ񹍉7��)�A�tz�S7�-Y820�H�<�J�7B��E�"Mɻtt�3��B���}�8�g@EeŁ0v�n�n�H:��Fm�˜�'�>���V���IV&O�ک�Mf���c�_FSӚ
Ԡ¨��*�/��gb3XE��1��or�%n�|�N�}uB�tlpO%zze����e\Zv��c¢�Q�F��}b�-˛����/J�KP���<�Z�bʱ�U8�(yس�Ȇ���2�(N��r<7C9�:#�O�Pk`�iۺ�B�,W4<=hl�X�ƌ|q�$�_�蜠�jz7���"���}�'� �j"���@�x:�M,6���B�p�����x��7ݯ�>�e��,:�����`%�.��+�ϺR(���4l9-��<̝������5U�52��~�%(�t���r��|b���ee_����R�F�^�{�?��:��ğ=Gˍ|��d軤��?�Ң_I+�·
Bc-uy���
y���L����;츜 [�6���t|�էm�B�;�83p3��F�c����q-���|� ��py鰜=J���'L�!���A]����ևv�*�Uyaj�@�Y��i6C� 0�,�hKL^��-�z�,���j{�Ͽ?:�l=s/�<ڷ�G��z�T3�)��Z����{	���W�>�W�/�T�s#A4�N&�tB>�z&�O4��h���{K��! �Ԕ���Fb>�1�^1x��5�`g�F��ܺ�MO]y��K0.{ƫ��q3(X�d#�f<[���W<Sd��02�J5.dO�7�}�#������'N�.���5��"�:���A��0��3
��^;��@���A���I�����ݹ1y=�k�j`�R]��>�ΥT�����g�F��=(,~�0U��fX̅�|
��7O��tԠVM�:��"�������Kr��M�w�]��IW�["���)�~!��)���bP��ɓK�.���6 lJO�����CF���N�`�QĕD�_�x>�����8�B%g�	�q�Su�V�?�@5��\8P��7ݴ`��l� v�2�osw�UD7k���9�n��ÙE�Ȱ���@`:��|uBDK(T8)Ű>T�oD@^��}�vut�T�e
([,�����bj@�m'�z_+��D����	��x�i��L�}���%bl�d�JZ��鼹���b���By�ZRE����	{Cꇻ)�/	����2AM(�{�'o��/^��2SS`d�)�e27��Z�i�7�h���7��c�p�qG�0��y��B�]�P
��Ƃ\I�ڕ�K�������
"��[�
�a�q�jߊ^���\bN��w�r>/��<�����kK��K(�i #�xН�Vb�4"�/@ٯ���6���6����GA��Ý�3��7�:`ɤ�	��Cu�V��*Бͽ�E���nsKXx�L�
׶��H�_[һ/��}�H/�V��ܘժ�$���Q CY �d"�piʘ����o��o�qIof+?�K?��p.M9���$:��!}xQ\�J��jt�[|ę�%�V��j�携B�pt�*�~ɒ2$��,P.|�tD�C�a9��aȖ�u�PI2d��w���c���B?��$��:~Z�@��-*��x�]z��_RV���Vb#��UC���KB�.u)g-��`�)��6��J"�pI$[�����d�9����
:���<*q��i��̡�h�����y2/�)IxyA�����,��B�g50��	����6�����bi^����sZ3�_�Y��-a"�$#Ȯ
upX<�*����N��rʡ��| 0��	�c�j����"������ONK�]\�"t���]wQ����]�T���P�)����;@6*�b����L����"�]���$]�,�ES<���9����"�,�}w�)�����ڢ|��X�&��4�l���G��Z��&ek��)t|�I���X,�V6��mF*f��>�z#�;ʸsøpD�&)�W��#����>r}�Q)�n�%9nFސ���R���]JUѲw)1C7Jn�)��������(U9P��e��>o��NW�便�d!(�d��L����N�HE2���  N�(�M&-(өl{Ʒ�g"�C�3Ϝ[��{�� �/�����h|��V{ܵ�NT1����kC*��h�pQ�be��7O��V��f6=�a7��iё�K�GL���n;}�r�ϝ���3Mk<	�O�����[�ՙA7tH�;
ɟ|�z��na��L��������j�Ja�:��6��9!>Y�[����^!�e�8\��[*�>K"�H���v����qQ���+�j���B�}
�����6��~�F!4�Mu���.����E� VcX�����3n��ԗX�M��^li��Ibs�{����s�Y��X�)@Rn�̭���Z#�3�?��EE�P~������Re��N�������n�4��
�È��2�nNO�Fc§���Ge���˼q�)�y���]X)y��] {{�$j� �*���I��BP���M"t}����R�m��rj%�Q�g��c���*��n�S`42S���-O�R~���z��I��6���5�h�Ŧtf�����t��Gv�4�?T�����U���M�9s��젩��!ß��?��V�l3}��\~W�8�\e�һ��4�o%����xC+����$ߗc�T')p^ɘ�AsR����v�Aw������}t#n��ƭ���V���&>jL�_޽,P��p�J6����I6��$?�[���HI��*�EA�V�Z�����'	�>��F��G����^����?vἈ`�*K����-W�}�
H*���r�E��`�_�sї�I�I  X_Ms۫BV�HG[7���K�0�� ��U��co��T���p��1��zd���c2��@�i�z@_m2�Ua_hA@����HE��Tka�R�Υ+ZיІ��?0l{���q"�jv�'�
�]ҍz�#����m�E��n4m�p*Qr�In%P�x(8���Ex��(��*i�+�&dG��+d�Ht<��#۞s��H:`��yN�G�$��pEG�O�Lf
gqDS=.��YLn#n6r$X�����D������]T|o� z�0�%a��<����g=��HyO�6?��j�X�lMr�A��b8�ߗQY�9�;�]?+�*��X��6�(:�6y>q�t� ��ReF��[������
��j��`=���W�KW!�Ҽ�/�|�7c+Q\�̘��=m�s����ȱx[N^��e��&�����X0Ɲ��EnUyGj����Z��s|�	~����s@���E��W���+9���@�z�1F��20X�,+�� ��es1}ނ�s@D��Qx`i�{�'���R���kY9��Θ��񫃂c�+��E8��L�&���YD�GU_(ӟY�WQ)�3��5�w�� �?I�?�!�x�g+S��W;7M�:Z OD�$�\��,�
��9(ց�,]D=�bS1z�T�d)KU�x�֏��=�\�vAkY�$��<���ύ9	6��pW�T�����ۮ�����+\�G�[��U<�'�
۸��<���"(|�g���4���Ks^1�
B��J�W�x���Դ�F�>��fO�qM$�Zª���vk`�������8h&�z��U�I�>��׹��B������{���LP�� ��k����yȕA�6�5�1�׮���n0�Fy�V��'TeA�%�Z�E���x��9�H��f+���z�Қ��G��#�{�,Eԓ[�'����I�F�q=9 �c9Y��~n=�F��@�\��.Z',����M�a�T�j~ L��z�10Ё�B$�?`@����*#�!9�1%j-!M�5\�v׋:Ɯg�ſ&x��^ii/�$YO��#G��TL�M'�͞_��f���wrv^sk# �₨�n�;���n����&3��{�[E�4`?g���|�Q�%����i���(~N�YrV�Yyf��ea!gzR��l�0���aS�]x�Ȕ8m.;*��Ѱ�G�e\IEźJc�h+�0����`rq҅RlB�Q�e���Z����!֝á��P����n�;Ba���ײU�Ƶd�5W�!����%�����r,�te�������>��l^���X�7�m�W�@7��wA�zl7D��%H�Zt����ò�
�An+��1	8�z���4�X�!l�r�-% ��G��P3�O�ܫ�ҷ*O�� $u�$p���2��u 5��F{�������ؾ/I�=H~	n�Vgݓ�u��+����c*x2��~f�����l��!�?xr�6�#��a����&0�և�?�µ�:	�򘫯kr-h�Qw�(�W����-[�=�/�v\� ��" �zQw�ӾP��F2��Ө�;�Q��0�e(߂�W�������>$�|E�X14�+)d*�<g�h
�(9����n���
x�
X�%n�%U#��+�� l�
���r*{�����_2�����6%W�d�D:ז���|
��d�LA��Vd���ĒW�g���H%g�T����v4ͥѓ�<����@�v����#�(�ܪ)�n�
�B�9w#(<�E�P|K�B�j(��=`I�f�G<w�-����9�+�FI'����y�(j�������?+z����g@�K A�����~>ueJ����7�<� �hP�)w�j�����&]��
	[a9$��B�ݥ8ǂ���Z���>���`����]7��jr�N��,����!���</�~������HCQy�5�,����DC]�`��A���(�<
�����_�&���u�	)C	?�<�pj6�T?hs���0s�)pȰ��.����O=I.Iu��Zʇ�u ��4��[�f:�?��++I���B�~���i!IG��=8�3%<L�]��U�M�N)�S����Z�\�2��� ;�,�K4��O�rI�d�cx/�v�v#"�ԕH����C0|R�ٍ��������V>�p�u�mg/���~ ���,٢��p~���H�x/��}�x��s���睗WQH�Ǣg�{�Ce�u��@�E�PW�s0�k���g��{�칣�)�w�|��L'�6�#,bI��6m��p2^F#u8A����������ҡ���3�g��N��N+@B�K�LsLKJ�=�7{�#��0�wO��r~���!��q�*��=~���xB	@�B�c$eR[�.�������Ľ5�ݯ;@�ao�i�m��پ��)�sghw��"�3�j�{A��>�Ux�������M��|�Z�Gp5��fK��Wr� f9���vв���X�]L��}�<c��SxF������iH�Ñ�V�<�,KH{$��r7ka+T��mP��� }�LD��V
(Q����#�����[���X�1�4&el�ͷ�i�В���ŕ)wH��:���!�������ԏ�R�����a9�	��)EY�R�� 3�i���ő ���u�UeW㪕��X������ ���)�ػ�$Px8d�`4?�V�늶�}B=<�GY*Ps^����:'b��P��%���踜J�R���n��a���c��4U�nv׋�P����CC4t[BM�eX�,1�oH��吏w�������¡	�����Xb0b=%ԭ|�r�dP:���w.�*z�ÔyR��ۥ�C�L��z'���8g��-�d�U�Ɂ�\w�'�9me�#�ow��gٝ��p���B^3sy�J���@��]�0�3�^7J�/<�Ė�{�~�hw���7����O�eb���~�T�·Q��o�����yK��jң�a�DL��e3�]�X`c���ݟT���[��N�?��� +��yG�4���x��H}�|�~�`��>�B��, ���%�ti��&I�������䝇n�ܼe��c��"JL
@|_;�C�Q�´?`d���4��c�닇���!B�oս[3��8t���ݡr����ˏjߩc��N'�̲�(~���4b�^N�V<�jd���~�ݘ��g����S|yO�)@(K����S��?` ����0U[o߃h]����~��^���yǶ&t�]�*Q59�ˣ�<�$K� ��o��o�_��$T�a�v:Z���N�>�; x�U�en��I1A{�!k:�FԨ��3���z�4Aqq��/��]ʌ��74o��}3�'䴪8��i�`���@&��BGl���ބ���AAkfS�:	<�`�O6iT#`w���L7� �77���r���N�	I��BL��s�wu)�D�QT�h]3EK"�8�XH�:�j#(JF�D��rP�+%#���܎-��;�m���+�8!~�����`@�h,mh�ۮ��� $�63��4�
��9���dZ�vLH�6�$b����Y�t>�螇�u�w���e�W���/��!GhZ�+4���t� �eo8 ��~Ѓ��Q�����8-��	�:N�S�Y�N�sͺ���j`L�[ƿ�,2r����`q��/�����a'��;gPƼ�bR������4��!�ob�p�p�UygZ�<n(�"8�[IRп���"�I�6M��c��>��Yř� ؗ�(n6IxǊm��M�{�tc�$�2���F�r)|Y��9;D!ȩY�S�B��T~~�p[�
����w�*����l�� ���?���R݆�����wp�w�sc�(5�g}#�����LI[j2�(J�sK���E�A�-]�V �#�o�8vL��$r�p�F��/>n���n�Z�Λ͏���=���;�Y���{�%z��~#���|�#�g���5혆( nL°���~\��J���B�#A�pfݜ��<p��z�M`e���x��f��e!?ĩ{$�ۿ��K�?W�D�� �5c�"�MM�:��g͎+�c�ߠKK!�(�y�n�f�,?�ԙe.H�]	q�6:���Z�4����8L�؇'����W��a[��j�v	?
C����$�3A�o���1<�m(�w�G�2�Д�q`�ѵ��x��8��3� v��3�"@�
�� 3�$&��B��l�P����p
��Ã���m�o�V�1�+�:��j�m��멚<��v%�ǩ�����n����r�M];�ƅ�C�.��=eLqA���1I/Q�ubk@b���j�`� � 81����H�L��o�DH�D������皔 ��
32t:�)S]�z�e>�V��~�|@&T?�9�p�v��}0�\�@�7���b��(ge����ir�^���|�?c���-����*�|\�[N'@z3���d��S�-�t����"�3�����|�'��X�<*�_�_Yi�+�&Epy��:B�u&aP��m��\.�*���M��g��:�X�73g2�`�c/pnr�Yʉ�}�,���3x:rS�y��� /X�*p�L���8��^��\ ޙ�T����䂺{�i�A*�ur��9�*��
������|�sh����E�����8q,����	g��w�<�TBӽ�h �T����,�ڽ���Y�������Д���Li��"�w�$:��6�I���
+�L�*�dv��H�S4s��}e9�+H��sr�^���U��/���*s�7l�HU����
�O`�v>UR�����Z��F��&"�:B�*	.�1���q��jYD ��RC��K�J#H��S� �6��D�f��r��;�If0/*pf��7~��8��#���� �XY�SA�Ψ�G�WQ�K�[�;�9�I9� ��4֑*�-u���+n�+X������u�.��W}�Q!�vEO�.�ˏ����5|�̂��۟�n6jS���M`���A�,��_�ۅ=���g�=F��&V����7A���OePT�'Rv[1tܔ;X=��13Uh~�U��ԝzc��
X�i����P-[�J��ެ��̎�B#�S�E�m�[>��IGs���n
 ��/�B�N�������rh/����5U@���c�0>f�,'��**HD�U0������C���7�m��ۊ��B��H��P+�D1q]���CBW3he�����9fF���a��Z&���XP�w�_�X*ef�
6"�x��'
��ڭ=0��!�da����g��B���ӆ�M�@pB��U��Z]3�d�bt�b�����&���s�\�?������2�Y��Q_z~���"Mѝ|�;�_�lK�!K�{�A������ �2���M�ܶ�;�i�ةҁQWnr�M���>[*�EK��8�:-��ZP	�3Q�W*�\����.t��g	����8���X�lG�z͊o�80�/��+�Du$�F2�G�e�Z�$�s��c�O���a�����dU˶�-�m����\i,��s�?�?��U���(����;,!dzdUϳ;�[���ny�y*l?ً��$"W���Fj�:X��^��al�o�-��Y"-U"�T��Wx��d�A�Y�)����<�[��.��/��ukx�q����))7�dU���7���-�}f�^�.Q� ZC��8����Y�`I���x�j>���>�0�}�-�)�����߱`OOzL���B:1����K��Cp=���d��rzzK���b�?7}q�]ɱS�_,%f�&�b�z�)f/��9(<Īv��_�z�"0��`~���d�3���Yd�;,�Np-:>�[���k
(�[��T)��� #�.?��ݫS0G�R%�d������Cg�^��f3{��� ��
vt�SK��T��!�-�����z�_�NG�]Vl�vAbTo�\b�{�h��Lp�T*]��"}�)xyF?O��[ۑ��>4h�I5#��i�C�\p��ɍ|�����$p�<e��D����k�����<t8A�}�R����6���g��(K	;]|]T���Vبsl���/��68���
��4�Qg�)e}�AQ�W]7Vۭ��IW���[vV���Ũ�XP=��B���zw=#H�H�qOo�܂��N?u�U ��C�����+AG,~�'<L���q80$UQm�q(�ҩ��E×�Aܒm�J6Gq/��ۗ�HQ5vo���Av@�����Qa�O�9��T�ԓ���h�)�	Zw'(�s.[fn�����p�hZ�7p4���6�y��L��j?���u����է�7�����;}�T�� F��O�Z����k���i�
���0�	�1;-��5D�y��������ORZ���O���5���h$Zż$�ң�㋳|�c���\>W���[�i�2V��g�6C��������jv��U��Q{T� $������3Ɨ��_;P>�c3���4u7�%����~�qe�ԏ��������;@L����k�����������ˌ$�y&>���05=�N�'��+:X����iKʔ<�+�˻-؊��Ζ[���D� {��M|/�ZMk�3��%(@��=��لb�>�ܺTzɣ�� �Dq��MprT>}����s�я	�e���u\���<�L�VG�����He�mph{�)5Zm��d7���(���cZ,��`U��VK]�U�Q�G~Hj���Y,��SϪ�/�\��-�S��e���׶�c�����P	m[�X���4�m�3�F ���k�c�C��S���f�U֮I�͸2�66�SE�O��0��ڕ`�8,��'��0�E��Iw�6n��S�6OQ�u�+�9�Ɠ���ie��?��|���Oρ�'(�ߒ1�۳%X�O���hr��S�3��`6\����I>g��Uͧ���6������g09d~O��=S0ӭﶢA;�#���
X������ŭQ:�t����?��$��6r�-R���
`
�s~��G�͌Pw3���՗��Jw���Dw�US������N4��������:B� �_�13���4�u�g��,�r5T{���5l���|g��<�~��>�?x�/F�bT�	�|�b-���:�=YT�b^ge��A�Tn.��� ,S��l�P'[�*l�^dUY�t�@o�T�0�,�#��4_[�ѼW�a��}�b 9�[2akY�#Dtϼq�	o�]�&2�H�o���kZh���=^I����%�t1�8:���K�b(�[�ػ�r=���Q�SA����y��g}�Tf���[UY.'_�E�m��%�C_�`8����KVehD��u���֯�g�}ƌz{�aSA2���:X�MbWN�kI�&�7m����'��/Q4��]������2���5�W1�oU����>4�ߓ%���b���]���%���on��!��1O�,V�	�a���c;#e�� ��Zz|ZOX�`�d�.���hu(��log_hO��)us&I ���K��;�`�F6���j�%�2���Z�t-�R"������>�o$*Ə�H�����Џ4b6P
� ���]�%!'��f�p�����/bP�ː.ң��+�/��'&z�V�tT4/~� ��$N	z��"��3��)eȎ���mTD/��Uĭ�$rG�ٖz��f�lD7�ߤL�|~u���y���c���Q�R��udGٻa�i^A ��k�H�s�e�4e&���ٞW���Z��'�ɖ�PQ��w��8��N�ݦg�B���.|�=��]y���z�7Gc������?d^Cl�`A��D��Ӝx�C�X�>�f�� 㑠�P�J�*��3�U#�d��� ,���5�� ���t�o�����jΧ .~�����:zv��-��� Y������t|U�^��9�QsD⍳Yr�>�o���^u�m��PאK��BjL3�֤��I���W ����\|��I#�eY�i���[7�|u�+�Oc� ���xv\U^R˷�Rص.�����XE2�`pY�Ē.U[��V��D'Q��t �Њ��,˻.N�i���j1�B�2�;"�z��WBBV&DV`��^
�hߔ�U�}�=b�B�@�g%X"3?f������f*�̞�+B�`=�|�?�D�+(
�]���\�Kq
��)k������nQ�|��ֆ.�Ȑ[O��(@��`퍌NŵR�yys�|G���6�����4c�h�Kx!�vG�vz^f���o�MRf*�C�gTWA�G��y�����O}8y\��U�u��t�(�gR�	�pT�>U�j�����ST�5��r4�m�9O`�D>"���R ���ue{4!�,��>B$���^Y8I��(��:��6�QN�_��/��'w��i�˓�b�!�D�������p�s=�s�U�"�]�&��焉��}]5�uF]����Ֆ�U�cҶzi�K97n���a��� \��c�D����R�zs7�����N2�pf��*�T8���&��(�穯�Ǯ-��B]=�� 18SOcbA��[�[��8z೒/���#�v0S�Lz��_H�q�X�%zy��Z6�Xl��)XԻ3Z����D�54O��x��l9lR�"�;�A#�(
/r_�s(��C�;%�1ӷ�殣��ː���N�h�ud���'=�Wz]�Pgr�7ͅ�NOl���?�=��*�5l����q+�ř�a�I 2kV�^<�%JY�qa���O�U�L�"�4�bgA��0w�&��L��h�#J"3��f�̻kvN��$�bf��072�#[��Z_ʶujgv��/G��`4��l��Ǖ&i��`�Ҧ��g�����U��:�.j
��f����U,�C�1.j�L�ˎ*�@�B�ӽr�I�:�'2v� �o%��@/���Rr�M}��4�Z�3�Y���GV���/��C��;������rz�ڜ�X�~(�`��]��	�w;OR��Un���qx���,G>��5'��������d9���Wd4/�0�>61�[�$�����+Z�9x�<x׍��jD^h���b�`\a �-�rY�q�H����ܶ�a��o\y�Ж9���H(�Y��o|-��qU�p%N'IG���KN̶f�,?E��e�����(څ�S� Z�m��l�T�6��ZgEP��TC�E/?��1'��6̼r��3���8]���W��|�l�ʰ��@fL����D)j0���h���SϨ��8�~K�u%\�$��?(V�.�A\�TJ��/ Z���h����Z����"b�S�+��Lt����(���g�q�~��"ą�TC�%�N���rä?��,���A�8�Ic��B'4�� ���s����]�h��N}�ÿ��c�0�G������G^��v�pS��]Ͱ�r���i^E�7�=?Q�H���Q&�v�7�r��@�A�5�{�|w�j���	�VG<���Y{>�E�rʼ���h��K��X`��Nv:��eu���_`��E����\գǴ�_���yYKh�$'@�����1����ڣ�m�	d@��G�,��4��R��DP8��H�QŹ�����1c{�������\�Dگ.R�j75ّ`�,����|?��+.�܀y?K�����9�9�������Y�}^���ԅ�1r>ǈ����:�$ACM��/�4m-��7)�����p�)�(YY�ID��I
����hT>�F�c[���N�<��6f�W<c��X�w�%t%!�v=0.F�I�����?�ƷvAsO��:��w�,k�`y
�빭���;�=D��4�`6/��I6b\�l(�	O_�鲢st//K`\;�c|'�� ���}��5[��G��Sr�Aн�?#�p�m�`#���UAоB|u���
щ��IK���`<Ix;9w؍��		@��J?�/�K���<����0�,#��9��Q����7�8�CD��@�	����X|��v�$t�F^v\�0���Kɣ���/s��y,hz�8����-�P��� �;l<C�>4F|Kd;�4u$E3���5����ˮ���wq�m���̤���N>x�91lr���:�5H��`��Va\��gE� ��+��;�!��'Q�]�QGjQ���K,��-t�hT�x��M��Uu�������j���cnR�xO�۵2~�U+-;��:	W�	���)��Fe¤��f�H�ȵD)�N���D�1w���+��w�"��d-uPvs���L�Q�|jE��qW+Ʊ)57��3���� W^f��=t��f�"d��h �MMc	���̹�?�>B����5�39@ *��r��YAV�od�~�q�>Hy�X���5�708�ձ��%��7�J��Gz��%�A>ʒ��<��ye'_��M{\��is5gs˨�߀�◀�q�<�� ��*%R`ЦhR�	?�a:�꽊��'�G��'Iv�DX6������1�9�h�lMz��M��a��o�>H���K�{i�wϯz<A�������d&��=��+�O�H�a��w��Ы	&���3�D{\1�.�Pj�˯��	HI�vԯ3;���8�>C@�Z�y�W 8���!��6$�:����JaB�������,�9y�Rf�gյx�ry�,�J�ҍ�K�:�9���,�a�$��}����D��s��L3z0����I�4��<����f��k��#Yj�U��'3�$N�؁�x#\� �,��C"f��bSŕ�[ñ�P^ʲ&|���8��k���I��µ�F���Jep�����3�2�ں�	'���oi��~�D�7yț4!�U�)���ojm"����/��-���2����e��R�|�H��eğ��=�9k�z�)�o�Wz�����]��S��He[�V���n>$s���A����!�1�1�,�.g0Y	FO^M�.��x��Pq��I�V0����?�,��L������K�Ytc�ֺ(#�%�E>�n�Sc5b�,�{?�MiZ��+�ù� cIv�K:�����a[�Q�����<«��ڻ"�pK�.��+)��P�I�9z�\:aPu�;�tEF��E�k\Wh�;e����N��25w8"{xX��P�I$�?gq�b�F���Hqd#R�qf��9.v�8�&R}���^�z^4���� Tmt��k�n�A�4D�abl��1���@����
) �[������ӖPk�`=w_d��1e��W������WK��>�,J�Q8Wƃ�ڟ��YO����C�8�����9�؇I9u��UH�^�:�a����@�/ߺ�iZ�f�ό��;�|��"4�*L�^{�n���u��J���3���-�Sp�)�k*`=��]h��ɋ��Vw���`;�1�N�J��A�ۿ�����E�۾pX�J������f#jyT)�.���X�ܘ
/;v���i"���"��^��00���tB�'�H�ӂhI��!�s���z.O�a
��eH@����VD��6���~_ۮ0Wy��:�3���^m�y���|����7�� ��3�\'Td����~~*OI�F�=��.�\���ÃB�h���<�ߓz�����u��4�ቺ�-+��z5�·%���9���U�>iսUe���E�W{�\!E��2���UsM(=B�&JO��[A�m�H���E4
�g�z�u�����)1ӟпQ�zA�hJ���喞��@�4����\�"�ޘ�'��S�� �׹���PR⪿�-��*�4w�}d1ZA1nK���D�ǋ���z��$8�s��45������Tk��4�/��K��)�a��u�M�G�h���OID�E�����\�g@I��ףP�ޱ����c���~1f;?q�sb6��2Uv��v�q}���ÓD߾8� �L���aH.�
�e	D|f�C�*�n��!���w�8K���Kn�fQ+2���/�A!�g�&v�.�#�>�����@6�@H����.��(�:�qHް�["�m��1͚�v:��F'�3�ɡl4 y�I��e����X*-��.��c�c�ϺGъض�c��
-��שּׂéI��-�3���ѐ{ o��e�\�
� �wO�8�(�6�J�+�N�?PL�i��a#�����mj9�K�I���!�O1j5���t_�}�g����!� ?e Aja��f�?�7�_��l��ٳF&�v��D�3(g$��Z5W�G:F�������Ζ�?�&�����4�^Yc퇻���$��q9���v��Ph�䊥��]�³ ��:���\�2�)�ʴ�����6�C�U��Q��,B�&�Mgx�DXvTL��'V�s?)*��#X��S�� ��s̳��#"��w��yՁ<��;uQ�7{$eC��D)Pw���}yڭ�M������n��3��
[�MDp�ȥ�Ӧ�mB/Q��u-�@7@y��ڨV�b1r�v������=)ȁ �|�
�[~�DiP���{Kʱ��N�:�U������˝�g�#�)9�禩�/�>XzFd���d��Q�匁�_�����pg)�Z�1�x�,4.�7Z=K���l"|h �
�2�ړ�Z���[C�0P0�z�}�>/��{q ܰli��v�B��6���XS"%Ժ�����C�_��n���a,��=�̣�F.K;�����⓶��P��	G�r�ew"��Ю:!�A�Z�[��æ���d��Ih}m-����rЉ�7Ѡ�Mձެv���$��/|���\/���:iQ��Z�s�-Ѕ���ߙu����K ��4���Z�#?9P��#�� "B���p�n��[	bBGP�c�
r0�J��3�t�/���p�?2Z0$��sSfT��0��!��[c���FM��ƃ�驢��Q�E>��A��I�yQ�O5�Yji<��^�:\��0��P3�q�'Li3n���z����}Ȭ�ƈ���t~���8',��r��jBx��+l����{��ւ"��j�m�^2ߐ�u|�5�/�5�˾I)ц�A�/1�@�31`2\�����?���]���߬�J
>P�/JUPb`s�Y~W�����'��@|R/L�F�� �W]0�����҈� ÍАb�u�,��j�;�>�Q�,�^�������+��Y�S%rn����N��7@��/:�þ	��UL}����
 �U��x$+�H$K�U��-;>.MAK�y�oQ���Q|v5�KX�G`b��gEq��������{ģ�hn��K��[1ڀt?�JEpFh�`"�4
������HH�(��Ҧ�,R�H�6+�6,������%Ն0�a�L9A$��+'
а����KnG�f��<̻���HŃ�k��G�����|֝m�I���FL�=m	5�Z�W�[9K���r xt���~��qo�λ�A�T8 nJ0CqY1��j��"���F�X��������Fo�D /߸�mՙj�,	
��se��<�U���:T~����fˋ�\�Y��W�) s�'��ȹ�&Zc�*��ĴB�.%H�Φ���4'rD3"H�{�Pǌ�H�|�޶���;:ZH���\�'�>��m:�3�OI"Q%"#��xf<�,^ښ^��5�GS��-�Z˄��(� �WX�F�"/�S�P|n)���n����
A ��B#\~�y3�*��"��+C�$S�P@Q�����z�(ʐ�m��!'�M�D�«UL
\�B�{2:�vvl])!�g��r<��#�w�Ju�L��$�8���Ƶ%��Ħq�����~�����V����UW�Z�?�8�F��ʊ������X����G�1��Ԛ�Y��C�!�q�$�����og�p���ӝ�0W��L�xr�J �-]�r��*mbŘ�U����u�D2�R���.�]f��R<��;7��GXEC�C;e�~���5Bİ�r�{���gO�Μ���{�
��x�H��A���v~N���q?��{�k�xb���_̂<��A���T:�Mv��Q���+ǓH;����Z���y���2g>z����S��ȟ�s��筻�1�2Tjiў<!	�L�+�}M���p[��]�7��� ���Tȓ���Q�e�oY]��
5�ރ0
�2I<���=�al��A�.;9ː�8}���R�f�g�hr3S�h�$,��K�h<'E�
����>j:5��tyk�y�u���i��~���c�8����´��ĕ[���+��?���)�A�O������
��X-�)
�N!&�2��D�|'*�����AQ��r�E*~�@*�_�[� X��
�����2v?�5�I��.	ϫ���-��g*���~�y)p�	�����A �I"j��¶��F��u�%.��������Wa�tp�.����;�Ѭ���o��Rp*`0� ��B��?&d�?�mVht�b�B� �G�}��p58��E�8���8!8�*����}wۧ�����k�@I�yZ|��y6�����T�F�c�M���L6Kpj��Lv��
e��?6���gY�@�S�t�x�S�ݾ��ޒO�����>�qp�$ل2��O�˸��9�zM�#h
��3��%�{pAV}a�:����1H�WΪ��Q:�Y��TIĜ35�-:�S��R�Y�����QL��UHHD*Z��TS�:�����<��1�D�r�!��
��-f�p�P��uI�H������l�b���_l�y��MT��.̘�}�UTe���+�Q�Z���'�8|rJ��lH�{wl�H�8ƪ~�2[ �dc%��Ј_���~sJ�X��
�{�~t���@��o�'i8�����%}��S[��,E'M6y��ecG�:�_"�O\��Hux7������e<m�2�~��	����l?_[���q��C>2�Y���Hp�E�Y�_(��Ŋ�Ω��V������^�Uà`'ܺ�UU�~ܶ%��K��ݳ�'v.荭�F+)]��G���O@�A��eN
tb�+�k8yƯ�&����,$��8�.�d���Z{�x]�e���<�]�lu�H��^k�s&�X=�.�!�:_t�_k����I��阶�Ւ�`��49_�z��sa0����6�{��N6�� �Q8���{\<3��jc}�dآlк���ƨ�$J�0�x_3��D0���Uo��O�Tb|kv�։������7�&�j���b?1e�{Y��{�*f��µ�2����� ����8�(�hm�Ї�m�@��I��mays&>�0 q�̥$`2��ء��@�1�M�:�ˠ�'C��~	G5��x�0�s�>5�������q�/���5/�'�s���?��\-���|L�I���E��ǖ2p������N竺[�PpPs�\͏gh�RM�]�C}V�sD��a/��N3H)��,��$�'��q�S��E$nǳ0,MU��z���������Ԧt1���h����L���=<NN���\�.K��~������3��"K^�����Ӭ$>����R�7�5��Iͽ�N�y�����U+��+��랸ʉ��%���w��߻t���P�0��j��E6��Z��?����љ�X�F�Q�������%���u�h �,�65��wY�r���-�g����[�-3���H���^�m�3���
����"�^$��F�^���/)��/����s��$ݘ^���벚I����ϞkY᫢�	)w ��޾9k%��L7P|�s��Y��8I�k���=G^���� ƚ��4��(�,�cV�@+�ۖ��BI�'[U��Y3��&*&�����g��J����2Ua_�7��Ɏ�{#��{a/�'Y���h��r�Ľ��+����2:OH���Oϙ���ۿ�x�婉Ԣ���
9��)�����un��C��#����B�A��_���q�'����|f��{��^8[5��X䃡�k2�������-IV�h|=�$S���K.ٶ��?�y������>'�_�Hj��|����,��]����g�:W�WcP�3����:������L�!M�TL$;#F�Q"���}�>j��BF�ڍ}D�ʕ5H�-廳U>��]�0G+�����3�[<O����F���X�g��ܤ��&Ѝf��8�����J���% ?�(�Zg<`�H�V�Q��R�SKoMx�
�h�բ�\:�vk��� �
���f��<饭�6E�3~&�:����I<��D�.�(ַ���nn;Êɫ~��+b���ح2<��Gh/�ϑ�Q�`Z�B�"�W���_�i�hJ��@-kI}U��D�d��y���Jך/R�J��wN��+�~��_�Yn�"%sHi�!��5�M������V�5p�K!����ln� 	-N)�}@���t����ؓ
n�{~�i}w�����7����G!��|,Cܙ'����>7c��ЊT�^j䧛�3)\�=RC�P<.�8��^IYR� %���0�EG	�`�H�6���,�~�^����Ќ��PK�@�&~b�RTf�I���#vOw�YŖ���zkX�������X��m4�3tƮ:��:���2�Z%���*�iׄb��-sK"5�_��b�k��Ze����8Ĕ6X��ŔUVǄ( ��^Ĺ6�!ȝ8������Xu��x���8B���a��� ���x�&)d��0,���^�c̹��G]��W��2��wr��v�C�G�[�;`:��<��)ĥ���~x���8��I���\~�)��X޿�:�ݽ_�h��)Yo���"b� ��Q7�ލ�ryN��|��s{E�Z$!HS�ym�Y�y���;ZT����+6�2e���ޮ���Q8����D7�1��(�յHYfJ��ܛ�L}dl|<�����Oe����X"m�i����9�:4��[9��G�����K.�1@l�26#'���@�W�\n .�Ejm�e@n��Z%�r��� ���y k�pJ�.��	[�S�U�~�AvT��qm�a����45!>B�R����FF٥��j�����k$s4��<�3��jj��zC��7�j];EU��1�d^�eڵ�(:xS�����-�v�����xJ+-`�Ή�(�H2v�"��a��T�\�8�HM�vJ�����~lL�O7���^_2]nR��R�B��?��|�<��1a5(�����̬ΗWهus]�%aJ��zȐ�R�uq��A���v^�E�Y����L^rUeƩЈ-Ǹ#vG74��pÆ(C��'�?��u���"�є�ϳ�Ȼ�c����Y��j?O<O9���~��W�_I?��/�J�ް��(9�H��4@'�XV
bV1�1$���*�ǹ1��ڦ�*���-�u6�ޘ�v]b�Y�\o��ia � E�z���6�E*��}o{�@�(I��>9��ŷ�y7��R\X��	��w����*�����͞���Y d���Rr���7K�Zd~�ʃ _�˼�^�[���ro�d�kx������Ki���F2��K����']��Cm
��}�3<��Mg$��/��0}|��R�֔����?=������_�����i�_{zoEuG�sPc�2�Eu����E2�i߄1���JB'�هS��9["ֽ��8�vFZ��Q�_�����0�¦��� �Þ� ~���f�XR&����@Fi�yL'%��}����b"�B�d��o/}�4��O�B�ꛑ�����)��?]��[�E���E�BĴ������hZR���%{%y i��W^`Vf������I���BϹ��C���%��_�T"�*����-���G��G(�6Ӵp�j�z��J#�2h�6�m��:$�zy#ү�2�M��&IV�&�~M�E�	�Q�{s,� 	[J>Jꮀ��;�.�M2:r�`���A�
����A@߱�A� �M�����{��PtKB��2�T��n(�/��R&�Q����K�>�ּB|� �vD4}`�m�T�����6ݒ�N�S��/Td O.�����R�i��_ wKM�s4���{���@g�w�{�oݳj�BX�ʷ��>�D/�w��2@P�
tbI��6�N_�~�ߕ=d�/�~��_���)�j�k�$���*��Wr�'Um>�4y̵��V�q�	��[W]�0���3-!I�j;�O ���r����0D�8d?�_�D�9�A���関Q3��G���}v�vV�4%�
� t����G�q�i�}��n&��^��E �6��� �e�B��Ь/͆��$9�c�n=+�� r{uN}�i�~���8+����*���8�=���Amx�<s{k��р{T77g�����C�*C�K(�J�FZ� ����=:���.����}/�6(@�L}~��Y�ĿۺI�l���A���S �Fc�Z�(r��u�<Q���b�R��:��?�K��S�vcTD�<�����k��&	0�I������A�mr	1�F��(�����ʨ����y?� ��P�ݿ�Co�S̼I�ׁ����/$��]����U��da��'��aT<yc˃�ø:(�g͕V�����q#���HM�/�7�E�ք_l{����
�٨�]�400��ғ�� ����t1�E�b�J劼�7A�g����u�P�V�3>CL+�g��e(QIӺ��N3jj,Ǐi�AeXl⨥�d�l/2,� $�(�ڠ$�1)���D�;Z��r|��8�����؏ O�aJ�B�Y_�L�`!hɺ�(�)�A�e�s7c[�Y�>�斢��1I�*Y<�Y�^��	7��j��eR�A�!3O���٩S�~5�i������x��=�
�����?
�o\�"�&K�J�_-�
<I��o�����M�j��3�����@E�3 ���z�J����ͳ�W9��\J3���D��1� ����/]�#���l�� �¡�OqМa�3�m�����?�ҠЉ �)#�n�j���K�5O|�^�z�~�Ѷ����)�
:�ٟe�Olv��*�D��H\.��z��ǒ4��	.:����0���˅��4���F�rʱ�&��1)�o#�_�Аk�J�t�E��nM��>����6N����L'h�3|���$�18��k�;ө���{��n`5l4N �@�&���� [���l�j��
V9+dh6Ad¢�a�8O���Nާ=�aa�6 a�*��~�N��1�-�#��	�,���š��)j|���	Y�<>
[���q+���k 2ͮ�����M�SfM�71Lq�S��E��2ṅ�\n�Lg�Z��7�,�$��1�?:�PI&���
oɧ��UD�DZ���w��D�gd��]�.�U�?����VaJ@�MH)�sQ�RE����c���+��hϦf�E�tڂ���p\�߄��yJ�P㯍P��v�5>nlw�	K%��^g�28E%�
�t
 9a�مC���)ֵJ�h��;H@*k�UO�J�Q����p��
C��E[\R�M�7��ƛ�VAV��wނ�*}�q���q��җ]�����������$��Co�ֲ?������Z��Ĵ�3����PcB9/u��*
���і�����ٮ ���3e`��{��u���FQL����-ܪy�V ��[�s�^���zEb�b'�^מ��S��e]9�H�T��l�> ���͔+�Tߦ�^w�pYQ���|2VH����lY�lU������I}�i<Ho�P�;r����^��F^V/�^Ocu���\�V٪�7ե��4Ωq��
�P �������K��v���v�k#�$4�S�f]��u��*�3�*�kD�ܨ�����RT�Jc�g64�x�H����M�a/	�?����3j���(]6��A�~��C6��W�y��Qd���ǯ*�!�2帎JN����8r6e��F�k���r� P:T�	�� Gz�UAŐ];�a�9��n��G�D_W[���$�d�׬箚Ț�XAb����o;�]B�B�
�,>n��)Ug�b���8A˷�����a�&���x����<]`|Q1���'R��Pڑf�6��QL��w�G�4�I����Y*Dye�>d��wz)]��Y"6��DH�BIP`C�N��W-![������F��Ò7D�u��M�I�8'���޻��M�
q����wӚ?Y�l%�k(�y���l����koȇ�@����=/�����l�r�U/��F�tj����T�0~D z�I���nF�A�������(ҿ�T�=���������̐aڗ�Ѐpm�^��yu��Oǌm��`�������`����Մ����� U�r���UU�*�u�kjt�={'��T�n_�1/y�B��f���ɍJM�\a�R����bT�l��qH��0q?r祼�r���M�ՒVCL��k�?q��B�?L����O[��]`��O�/���@K���k��`9���C6z@��^����?SN)���q�_�(�1v��8ˬ�*������,G�E�,���gr�F�3���C-�Ab_J�v�<��Hk֗`ZO���p��t���5.w�ݵ4���õe�����5@gf�6.&I�o�w��_��8��{q�~��M�f�J#)=�d�/e_�!���q�̰����ssf�!R �:K�rm��B0"s��Wt����ZM��%�6�;�J��D��p��$���r�/��a*DNFG��e��֢����'Ϫ7\����q�bgA�!���9�E�݃�.^��C�4a� %$�]��"v�4�Y�Xo-������A�8Xg�:���4�������*���6�߭�����捼%�Y#V3�V�7�,�19���x��tuh$�.�#x��=?Ƅ5z���J�&���+?zI���|܁z#�:�p�[�6�PSU���P��B��Vt>&���Q�|"��bhI�<a�y�bUm�����d�i0�}s�\%�b_W�Gfs��գ2��A�X3�g
6�=�3���Z�]	E��o�u�Z���8��__���OX����TQK��%ʳ$��xf���I��&K�c�vϜ� �(������L1d�Ux"X��f�I�*�S�����cK�8�6�gC��~w�fS��E��u����9�OQT^@4w���IL-25ߥ_K��x��	��.R�#ƕ���)���ji�����Bq����� ��N5��sH/�!Vo��YR�+M���j���Or6�3�i{ԧ�H��ґδ��c�Yԯ���O{8| dp$�����E#Z�c�?� N̻�e�c����Rҥ1,�!`�:-�.��C��OŪ��C��_N���O��|s%JNC̬47oz0>�-c0281y���ʤc�id��ţ��]�j�E*3]�ҟpLx���7�;�sm5޺ٗ+i�j�O�AT�A�PaĽ�?��>�P�.�d��yaaD�%����f��B��2
ä́h�8ԔdW�і����
���7�W�x��)���~���*C-��OXΤ�n�T����0<P���;���ക�yF�1�UT,���Ĕ�Js�-�����mJ�<>�e�r�4�r�cm��5t��č�Ј�&`�~���o��h��]i�1�&o�%�l��F�X{^6Ca稚��|��/��vZ��.�[9��N����J�?L�-���.�i�]ޤ�2��b�h��*�8+/8~�HY��j��v��4l��2m��H�R��p�:�`}���f���l�Pde���9�l�����4�, ���d��(�z`�ę�q(>w�>sY������q}�>���c��?A����t}�d����E@�(��e��|~?�_���>EC�g�W�PEq�����Gz䙜5YX��DR�g�ݸ�u^Qjl[$�[�OZ���Y
iC>Ir�1qyVN"�ᗦ�m�4���Cο�r�]�I��F���5���*j�<6(�_��J�nt���}��w5|������d�a)i�%�'Jb��0QĜ�X��	���J$��2S�S\���Mq"�3ag�m�M�lc�js 2������4L)ٺ>�� �����l2���m�ل��N���8@
~o��)i0&2B���N����3�$�S��_��3�5޷�S�u�|�%����AD�cz�u���q5���NC@�8Jj�䝹|��O���20�{���:����zM��z9��M�_�`E�:��w�t)M�T𑉐��Mm��a�<�U^� O�]��ȇ��N��JTw>�by�J/f�Fh��������Q!���DRż�5�p����ǚA�6&�%�k��|�ү�fzU+kp��
ܙ�' lj3���"EzP&�A!�W8��Q��~Iq��3�XMȰ����i�^���� ��s���4��1���n�pNɴ���_�xgj������7��<�?����k8�Pb�i�4�/L-���sR��[��=k�P�Ĝ��7C�5�?4�hΚ���͑7�]g�li����#�[��aS}����i,79÷����T���~�eJ;B;�<���P%�D;���	�Y�ߥ.?����BM����*���;�P�����/
�y�7��b'
F�4��aƅ�:�v�v�1�jOVA��u�K���	dQ܁˟�ǹ��Α��J���%�g���Q�[\P
�3�Q�t��9+<2N�z��S��e����H(+�	�����'+ �$m���B&��h������.�%�Z������'S��Ǒ���A\$��
��I4�km0 ��>v�!L k� x�Q@�^�#gS.�ܯPʀ5@K�tj`�Y�(�陾п0\E�8����*�O6��b,ik�&ao���1U����A��Qqㇸ&�k����x	޲�Jn�qMm펢zߙ�f>��:%�C �d���7����u"=J��d�����`P%��+VQES��<�]�WAL}s��,�+س��)��6|�>ʑ+5�M9_,��!X�}�����؎)�������U��.��ֻfT�>MP�#������E{�����������gy�=Mک�מy��Z��S"R;��l!4s��Deh ��\O_�������>�xJ�Evɠ-Ur�'�Z��@�󩄲x0s�,N�*&P,h@���d凰�~e�8�Mk?a��oyHD�Y�>�'Q��u���!�V���>ϝ��8��r ��x�5�\8�5(O�)	���X�og�p��d�3Ta0�(pb_)�P�l��	���Y�i���{��~��L�Į����`�� ;e�9�w�0��f8�dgiuX ��*�ƇiݨY��d4�`�Ň�p�2jD�dN����
���wh����H�eK��^�����R2�t�a� �ِ�49�4Ď�Mty��7�_���
{'!�����=iu������.n����ѳ^�7ϵ���8]��R�f m9����S$��ւ���b`=M��:2S� ��Og�]2�b�N���Be������r]+D9>ə*[ |ҵ��F5t��Ӷ��n
*8k`�
��6�������(�p4�s���\oЉ4�<���W��K��큔#��jI��D}��Vغ�������84�/���вN���m�D�����M/MY֌�f�KBx!���͏`��#�s;�ׁ5��K����6�u'W�O��[E"����Tei��EK�JS����`R�$�U[;y�Z�>	��Y��<S������c���lT��9�̡&���4���":=W�^������.��9<8$�JoJWfn�ij ~bV-�A� ���(@�h.Yw1��t�\%g��Őx���(?R#���z]M�V^9�g��ȱ��o܈�e��oEݕXE2��7�^���k�"�Z=7��$2�i���p�p���*P�
U���������bțB�NF>�{"��ޓ4\�q�vB�Gx6yF���:�5�� �`i�m��C}������x�����V`������f@ܕ�wx��)R�������	w�Ϟ�P̬+aQɩN�E{b=��+c�6�V��	�N��J>�����V��k� w,��<�q�+^�>��2D'/�:�����(:�u�0U	ɠ�7�4`��H�O%@`a)�kW���x���O�ǖ�A�����ۙ����u��ckZʜ�3������Z��K����z/L�t����	�J��iRK�>�+�@_���j��iZW��#���n׬O�|`���#Y�}�/��"���ϻq�u�B`e��_�X���bv�����'�/_W���g�����c�ϴy���;����f��`�:Fm�����Je0$L:X��%1Hf���&g���eT<؃��a�@�So�/�0�?�O�'�+Z����*!H��U�?��U�;���<��Nl�`wT�����)~�\�,�H�	�--�Kf����.�:�Xe%3�𻺻��/I����/!u
�AP3dy�sGL��t�w��O���c%�D�(ٞԾywr��U��ɥ��YS9������K��}����k�S�T�}*�6(�jr��˱9�������F��wR2��A�qd6�3�H��F9j���Ү#�3�4.z��='uE� ;�Y3�-ft�6ε�=.RBR�s�@v�̇B���Z"�;P-$O{@�y)#�"��$M�3O�P��܀��G�c�D��q߬������m�uؐ�`0+h�\�;�EZ�P1��T1�`�M!-��_ɀm���ҽpqi���e!j|�-*]a� �^Hp�P/h!UoJiL���"�n��_�!#I�k.��٥?��?���е�Gb+�wO�cAe8��3+�-����R-���Sr��!&Ժ%7����{T?�dGQG���2�(�g	�m����n����%p���u�ɦ��9rxM��0��6!M��:���ub���>�dn��N�RpB`�u�o�Z�_Εq�Vg��w���;6w :�3.�VfaX �8/4ڂ!o5Lr��~��ñ5vu�̭����-x�ԛ�B��*qX��W R��L�@3��uMW#�\�������3��7���P�B�x��K���:��ũ���j�Ŀ��	�ak=��N�����v�ij�Q��**crh�tð}�v�V�'mwf�Q����Ԧ�N��ڊ����
���30�&���ham��Hrև����1JU0ٲ�q���i�8v�_.��+��~��W3z&��	'�[?�O�h���F�Q*�ĩ�Η�pt뢔�a�SI~�/R	�Tq��5���y;��uF���_����i-�p�N�dkL��v\�}*	 xk��g0}<�$�M�-�˕��V$�b��^�J8��[Hο�Sb�P�0h�.�t�`�VW}{+ FT{5S��{HC��X{5g���z�-�fjne{���.�,l+�5�3;l]?�/?ynW� ��s��]�:v�k���,=0%
4�Ӊe�m5�(�|뷄�pb�ӶZj��w����۪��@�����X��o�֯��/F�`�}6�����BG�a��ձ�T�"�m��R�=����4}��Lo�6�w��r`tS��v��bX������Z��������I��W����=�i�� �k�eh�2��z��*����b��S��ҥ�Y�c��JuK ����F|�Hy�z�iO������֬-�}ضR�]�>9��9D�t" �ga�g\��l��VtD��Hm�ܳ�+�&�]蚤��ת�ܦ?Ҁ�E�k��~4q���v��
x���ʟ�����Ri�ν�FY����_�l��!?B��K�� MT<O�R���$�:p
�/U�yg�i]?��[ тߌ^�Y�d�|y
�6]��/V]������m���i���E>�단���@,�m���x��dV�e�͜��6�>2��mUkJ+�U~���4k�A]_8~�ڻso( $X�Ѝhj�hV���g�n�nV��T㺙��:].���Y�R`��^}Wy�q �ê(۷�;�V�W��P%`��' {��S�a��2&s���I�RXy�Ønm�o44���%&'䯫߉�֟TRz����{� ��D2�X*>4���hq1�l@'D"u��j�0��ɧ���P¬���:G�ǿ�j��X0�7or1++]��$��HZ"����~K"��?l��@}LQw5��� ���b�d��v6ZZ_r����k�Cﬣ�@�?����(Eq��,Mi���2�}�������VW��\+�u���E��̱�����&I�D�(�:EH�l�t0Nk��nc ��<j�7�w�3��[+~�\��x۞��4p������ɭ���u�nTNK啂��?�#-������\a����%�t&�TA ag��U!�>ZB��h˙���~�کzv����:v����#�gP����%|/�42��5��	�mY�떦n�-�<��piY=��:��Gw�������N�O�����:�$���&.8<�A�J����E��%H��xR�LG�6S����LC-BN�P�0%���	���Ξji�]�Ký��~�?j��&�3u���>j�b��/�r���?Q�	<�.�ZH�/9��F�T5]-7U's�a-�����ꢪ0��3�̺��n~ƃ�Gə�����mmآk})�:7���9i�_�6���� c���Y@�b��S���{�OM�h�j^#�n�J��H �+�k�����-�X	_Xi�Z��Dtw���m	� p'�f8O����O�+���?�"~ {�hr�*�Lg�V�!�TS��C�&n�ˉ,Q��X	�W~,U�Z��bioL�Ň;P�ȩ��V��;G��3O���BRnL���Է�D����ҊW�&ϳJ�&�ޝp������d&���[A�7�˲U���&m�lS$�υ��� +��a`Az/��v���z���!X
�����6�TS�n��(l[t7�b��R:��}�)o��=~���6�L�'��Zg$8[{�T�#�	Ib-^��� >�����qf�<�Ly8�q�*rx��O��Փl��.t��=A3�,��D�a�*tr� =���+	Q���u�z�D�+�i�_�K�vh�"��mzԯ�k��Wyy%,��JV�V ��~2~u=�w9\^($CRa6WDpzY1�-i�a�~#yWp
߰�mIu���q@�h��b��m�eQ������<x�����{�JR��q�Y��Z3�Q�6���3鵒!�	���p���혓��䕲X�p�i���Z0av[�bHd�R�朱<��\�U�9G ���z��	Q��?��`��SfT��h�x1���k\V���;Q�����U�����c�=�Aǀ�2��q�xo(���,o\�f��4
U�b1�&��ȋΫ���:��
J8�y���[��TĘ�;�֜�q�\�f�x�Ո9�I��!��w�TZ6���&����K΢Jn�+��S��"
�O�$�� 䒵��_)I��5�c�����@��tZ��-4�O��}Q#"l�Ԫ��罏nW���4�[�*A	B�T�7I%vQ���-\؈�j�I)�k=%>8������M�XG��	�=ﲫ[�Ñ6n�#
��>HE
)�Ά
��-���d���)8�`��#��g���&�w�g�>!��T���ƛ$�V�h��$"�,�¡�V\TJ�������s66QҲu��_L�H�%
�7�>F��&,|�"��5��S]:������F��E��9m��V�D0$ ��l4�<J�Pz��k^��ysm�4{��@�yJ33mL�9�O� �_1�&�'��B��S��K�]-W���9�=,�r��L�)�FG�� �}c��]��S^���q�o,����i�?��{�{�����LnA��A{�|�l��J��h��Z@AT�p��k��^m5uV��l@������)y+?�����B�΁���ɤ���g�w~�!�xˉ�m��XF;�/�.~Y���!��.�۫�>��-������Zǚ��?�(.kW��`���u�&�ԾubG�2��W��8�/���G��d4r��l{�b��|��+�p�m\�h���r��!W#�YC��{�@Rn��&��;��qy����c$��>Y����nh�^���Bט�����4�(Ӹ=�����b#!�X��6��!a���F�p��/I�b�wW��������uw�r���V
n.���^������S���hQm�ӷ	�^&P����^����=x��2,a!C� �Dp�J�NAp�c�Y��X��jh�W�n

�lMفև�_q����:P��<w���S�P��W�'��W���聶�N�����Y����Ě��'^��X�񆨢�7��pk G*>�Y���45'����m������y���i:�'|\�E�Lb�E�l*�",$<z�r�����J��>!jzv��%�BpD.��d��m'W�m�z~#�]�@b�Ù�����8�(����y"�Z�⹆���Y��⦈���,��b�-��jӋ��� ~��y8*��E��a�bJ�I2W��T�\�{	a��>��'���;���%�?���Xk|�Z�+k�D��Ze��s��@����\�����HtAΔV���n�$k���]��SH�>a��UA?���H�[�G_uԃ�ɪXr��C�1�ʫ�����"����Η�F
	�}F{}��qG�s�ha�:.�u��<���U&'�R�~�'O�Ѩm�O> X�l[m�R,��E!m��y7�(h��6�T�k���&U�������KU�&���/�\(oj�/�$dy�*����b.i/`��#���8�T���7��"it�&�2��X�ҍ��Cy�;���ˬ��E�eIRH�o��	��}�fӓsu0�7&�z7���Z,���HK��y�v}� }��bTPb��~�T�_8ZŒ��{Hl������k�ǩx\H$M��W���!jᏅw������TRBK3ZK��:& "+�����!�Q��hڹ�� v�T�A�J�J��۞Y���'��ֳTNo��A�'#�2��]z�����WQ��E�8,ߴN���f�}ĝ���s�ǚ�[�z��D���0:�N��F�`��9�"�P�,*UY�� ��q�?�����R� =0�� H�&ɴa��ue�Q�A��@Z�#���Q
�0g���U�
ͿE�⏅�V�Ǡ.l�?�*C�T�)������-iU�Xv>��7F���I�Q����,@D�VG�n�_��Q��ߦ���M��ܐu^SAV�S�:w?# ��
 �~+��&�����c�l e�	S ![c�ci�-1�>�ea
�1���T=䎠��o�Ox�np� 3�������@�	K�� �8�F��_g3�eh�d��~�l��J�����!�	,Z��L��N�2}���?�va±�6�G:|�#����r���kC�k�]#mv3� X{^�>%nnT7��C.�P�5�/��<r������Hy��N�N'�3�F�qq1Φ߇�sÞ��� �{N�ʢ�m�-H>ފ�jZԖu�m�������]��^��%��e�J����С0`8.1R��\��A�娞q�6��8�!�"��(h@Ũ�������*�[����w�j��sBXXzB�<�ݎz^a:pD�n"�O��,d�zBf���4h���!"T�օ@v�3�fy����˩�$������n*L�2	$f��8?�k��E�s��q�%.P����o�ǣ�C6h���ow�|�i�,E�h�)���i��K����xd�?H&�-�}H�l���O8�7�9���vJ!�6<#����0��\Q�)�ʐ�>",���h�kAc�]O��"G��3�}�i#X'+�k�P�]^�C�,���=R��i41���G$}�i���6��fl�=�o%C��V�`��G��� p�3;��T�N��ߋqȑRa��2�[^�@S'>y�B�����T�CM�	3�1�&��Buf�����#?�!L����a9 _"�L���Ѱ�j�r$�c@�,@�m}N��dr?�+�U���ݸ_f�׈�)���Zڮ���0R�g;��a�&؉:߰P��0Z�
�R_�0����}��ʙ��؟�B7�ut�F��q����g�к!�l�J�?�I�Pc*q�IP�� ���]��ܩ��i�ҭ�|�Km���lE����M+�q"��mO:�(����h�Z2"���ѽ�vʯ�U4N��5{Ae��I�G����F��G�g����N�� 5x���G�K�L�0"�J�)�Ƃ �
,H$N�����%L��q�E�&�.���	�fpnpblk�j��6Z�Q��3�b���!���M؍�u��̗xŮ-��/p�j>o��&�T(���/9�n\&(���~z�=�h�.S�V��q���Z���M�`s�@'Ȩ��0�^���p�Xm�8yP b�M��^����Z����� d��$���dײw��Ju������70���� �	Ü�u�>����Z%�xd��T�~�#SAe�Kf�c��.��,�f���:��)��û]���-B�_�	y�bb�7��d��b2c�����Bg�6Bӆ1��D����d��>dPܸfOb-���K���|��Ml�Y���L,�w)�dh�����+7�e94�Pc ��Na�P;FF0e�Ҙ��ĸ)�.ls��iidU���ژ��N!{��ژ-�r[?�P�_�V�V�>����ӥ&���O�H^$����������?��n��<��k���|ȿ�@���ũ�C�e��sa�^�i�-a��=n�J�B��7��7�;����΋B>d���'�R�$g��'jK)�0*�M��v�ؓb�kE��K�`��KY�9��1��1��.z+bX�E��lu�vi�c��EJ[L��*'�26�sy׼�ީ�j�T�� z*��=�g��=���s�A�PN�ăf�������k��6g��D���R~��=~jeɾ���Y�8HC {�|�q��?��X���-�Ai�������9�y���P�]��3#����+q�U\�s2x�����K��&͑���%a��o,�܍���;��a��R ��9�B��G�>�NL@�h�<3yƫw���7��5��w��6$dM�h*�d8����N$�F �����c�����
����X����*�\��1��y�ܔŻE��	���Q-F�u��~'�H���n|c���
;6N�g|�O�\0ú�@�B�_�q�#0������Ϣ��\��ec������u`�Xt���ES��V;Py[b�B~v�+�kzp2���BK0#�;VWl��j�xa>���"H��
%俛Ӎ e�_��d� *�%D��	ꨇ��~��B�zѪ��"�3�d������8�7"��O,׈?OM�3�b�Q�m�5�S�9%u�v?�8 \�U�����WO����$�`��|9�A���&�i�ކ��AH\�v��$�2lwh+�/�ǺI���<"Dӹb��v#�sӺj����HҨ��l�7:��m�����u��77V>:�d6��)�����ǵ�P��8F��T}H3lp�N�b�i�@2�ZiP���e��:N��w�e9N�YKl�2�"�<	�'�7?,+jи5(7�3����h#rf������֖��Ӡ>�H��s�L�K�;5+cY�}sk�aoT�QC�-�	<�"���+P푫����i�.hg	���>��@g�;�WG��_�(�����Zw{��b��f�g7Y�'Jb̹�s�Zw4����Q���05`����5���U�i�V}���� ����:��ՠ����nd�.@>#kL�4.�if<��*���^ƷHy�M�[�ܒ)�Ur�]�ç���D��ILr@lFsV�
� l֧����+�13���,��d���k��:���!�|��J���=��&�|w�w���>����0(��"�x��{EL�st��S�Zu3Ç3�p�}Ez��B?��%=��eq�������E�!�Վs��^ڛ	u��_i�:|
�� ���۟#�)�!҄T�X��˜�YT;R>�����Z�u�����\�kj�6�q~��&o�z���?=���2}�0�6�����ȑ�\1o�Q]_!j��\�<��c%��lv}W)���.�U�t�=��J�Ҏ�؀|���z�2YVI�,9�,Q�������d���1��A��K�2�#��~�'יn�a�5��zp����{�z2��"[be$h5鴴�i�D�(� ~~�V��,�4�<�B�E>���R�L�,�_..��kF&i��,2�S�{B�`\#�YJ�ڒ�b��-���%��޸�SK +a���Ľ�I�'��M +�TvM�훓��^M�����@)	��RZ6_>M@v��ŮUE��bg�A�ݘP����rJ�bÔ����]9�^�[�ґew	���;��{����t��Q�K����� �t-���~�wr(ku4��	b�-a���R�\jM�����Ujd��'����d���\���ͬ�$��nJTWG@S��{��rn���Pp�� i��@uVUT
�.K�U'3-��c�@�XJ��������j~=P!�����yuX����F�a�v<��#�h=p��2ig53R}��TL$�a1|��1��:��ɬ�AK@�?_���G�b�ׂӯ2��CP��Rn;����+j��
����3�Q�"��"(�EN�Zo-g-��A�Ǥ����h,��u��1�0�+�L�ؠ�t��4�Q6#Mo;��`&����vRm�r(�f��ʮ3��4&����1d=��F����P⨨l��v��s���ׯ  .!ߎ�O�竻|_CSˮ�/��ӪdY[�f!�tFa]ؑB�#[Mf���-�
X�֊�1�㮺%.8�^Wa����7p9�W����)b���$t��=3n,j�쉮=�Y�58���5� 6���!z]l�P��Қ��v�.l�x؍���;aHk��e�xX���jq�˔��0�>��*��9m=%�i|f*�D4�Ex?���)8��{���؆�y��<3�\��u��8�P(� bC�#�����@OX�����W�x�� �d�ֺ��w9��&}�g�#ps}�iH�ҡ���+l���ܕmm�r���q!��4�ѠC:�߱�R�sE�&�(H�
.#(�n�4�8�kD��՞���l~�����ΰg�y��@�o��4B9�����7�L����3��Kk(�"ȩd��r<��ea3������X����Xg��{�R�����@{)k�a��8fz:����-g������t�j��p�Td�J�(H0ON�U��6yZʾ5����YΊ��(�� ��Z�|�+�D����ax
29�>n_>��Ny/z��������|�I���^����T���b�Z�)"D2���*�'։��Z$��V�q*`^�|��Y�R_9�cl��o��ͨ	�_��N�i��m��A"Ǖ��`tp��[q�,��T՘��-O7���e˝�q�2���D����E�f�)73`�B!�b���?�:ɬ���,�111Y�Kw����m(#�o�`�������D�����a^G���x�]�o/G�<�������(�Gޢ*�Pú��s�0Q���+ڌ�Z%8B ��>�Zɜʌ!<�����&i�&,<�$fc'��|���MJq5��笩@l�!�-��'A��j�
�;��uo>�
�3ѿ��o��a��(��$��S6�Hrt�r���?�y1�+ß�x{��n��BZш�V�QcƂ�=��q�*Έ�W)p}	�)bq��k��[�M2�tډ���ꖢJ�[�:.���÷bN�[ӄT�k�/*��@Rӹ(���R��7��GC|�z` ����6��^�Q�X��b'�4����ߵD07:���fI�����J	�4������R���ʰ��Pm�ۢ�*��HQ���*���,x[z�D��?�������Õ�$�/�~2��Zߣ�9�Y����w����Xy��:�^W��w���6��j
	Q+�8%�*9�ڃ�~-=�hxD��Z2�c�Mt�Ȃ��K7�A0V�� -���ҿ>�"$5�c|�F�>|'X^I3P鵠I�(����E^N�X�7���pk�v�A9�H�sX�}�C]��=~8[��J+j�2M�'��#� 3��E�k+�.V���"��N/��Af���L����T�eݑ7B]����ajG T!����vl쁸3�a
Fbw������� �[�L|�<��T\`BD�d��3K�_8ԧ��+�NӤJ��[Ȉͯ!�$�E�����\�xn>J#��`D��ttZ}��!DW���0��]f�·7o{�a3��&ĩ��F}�pTZ���͉���NB˶֞;uF�1�7t�w��:5������.W;�Z����5�B��Uչ�1-�A����LJ����6*��-�*;3`�D�ڡ�W���^>?W�h�J�.���vc+p�@���_�W��ʎ.���2lNJ���vJf޽d�~����q�7��d�B�
��S&���=�!�И0C8���0�"r�R��r�E]ccՙ΋!/t ا:ߦ��r����ILf�炒Z�&��zx�fe`"�6���g��>��1�C�\ ƻ�@���+B�P�Շ�~z��c\}�C���UmI܏Ҍ8[`�ag5�3i��tg��j]�e�*f�C���G�/��S��;h�cc�����%*��Qz5E�8��:}%(�n�&Eȧ��J��:*�ђId��]׽o>��#]jJS4P�հ\�b:��&U.
X�N ���
@���� J��M�X'�+��N�(��x#Hs b�MV#�!�}ao�ͮ,Een�f�o9��i�Ϙ�_r�JR!��#p�c:�{���[���vK��~q��`!��j�7��5	�N՘.=�E�!��v�}{�p�O�"�J�w_���c9{�,D���P��x�O;. �I�,oou�u^Y�ˁk6�Z����A������^hhKp�v��;�7��|�<��q���2�O_���N�K��]4��[�1���=i�
Ը
�$�/����Cf��������gط9��;+�k+v��!�X��8���	�آ6���:�
yM�s��XR��:"��k�h7����A#��n�MlN\p�T}z�K݀�����r�c*7��A����9�w�?x&[�ׄ*�*���I�.cz��Ǘ5�o�������R��|���H�C�5QM����P���{9'a������^�l�V�k8�+n�S9���DRߵQB.�:d������9Y�N�;��b¿N�Iu�r9uY�<�?�:��G�}��l�P�Ej<�ۋ ,kל 6,̃i�������E8mZ�s�>;L/����1�3f=�5{��&�Z�h�����N�������Ӑz�FF�Ҭ����C��嶖
=��N�Eh�O��؄�ފ��d���3�o�E��̔�8�fj��b.�و���U8�a��
aG�lr��W+u��,�����\(|��f" ����$����H*��{�>r��3Ĩ�4�<�n�PyDEK(��P�hI����=�o�j�w���Q���`�sj�7��~��c����)~�.����j� �������a��I�k�Z8�eA`ko,\uQ7���y<L�x��t�z�CĶ����\�h��#�)s��j������MC!��o^¯�$W����
/Lx⚡�,���+�2��\�=�o�ުl������$�/dǚ$d�8�&I}�~�_�k@�0m��B�XC�l�笐�`�H�y�\o<�sf"�Ȟ�AO�9�){s�왽�I�	�ƚY�%�E���#A��_�s/���L�W��s����zP��뙪�dCP�p�L<ټ�g����o�)$&�՞�q��;gr}�;~�Y����a��� ���!H��O�C�j�6nF�W	�%_ػ��u1�׽ERj�>H�Y'�Ǘb��;�Nٍ�7�Հ����BQ��l���O��U*�dILP��݌�7�"G���z�XINȉ>!������V�����|�?�8��s~�|�F�Mz	d�+�("�ӑX�Z��EnS�jU��Ȱg�2���O"^h6�Wq��y�)"�'~T�.]E�a�5�z�K�xb��"��]�`y��S���˛���x�^V'�� ��.���\G'R�ŋU���3�{��C҆���Є� II���=�� ���06�O���96��z��c��E�� �!U��&"�@����M9\\ʫհ����7w���TЛ�W�>7;��d���z��δ�WԬ�di�q�ӹ��tR���D����cT� 4~U�:�LF���Q�	���j7kD�7�eg^dTֱG����
>��4'BN���o�'��u:c�&F�%���n>g�e��K*̞}����/�;jwk��`s��ר��]ДÉ��N8��,7]|�D��Z�(�kGE1ţ�Nusw�B�H���3l2UY�&��K[l��+�m���#�"�6�'x_� 96'��t&]����>�	__�����Q; t�,�"�b�c���|u M0���Pe(l�/��d��cBKtvō�m��s�\������Q�r�# ��փ��k7VYͼ�4�E�<��V(��^���f�����w�&��F#��S�	�vNE0k)��a���j��_%kq��e�6�� I"
��o4�JC�Ö���X�������_�� 8gפM�v}W `�gv�� /������:\ժ�����
5��G���cVa��M�U"�u��@����Rν�R�xU� ��u�-~e��:cF>J�t'&��[YƍJk��u&�y;;�v17�׈�������P�k�}l��8rp �B�����af
L�8�uz�?��4��$\�7�S�@�y��_5�y��x>d*�
��	X�)����ze �Z�}i��ֲP�EV�(*~�om�[���+C5��r��h(p��j��T��M R���Z�HG׬����������*�!�͸�F��^:�m�G���g90G/�3�_ v�c/S$�J�
X�����	v�Xg/�8e�a��#�n]�l��я=�[��`�i�����X��j`<�Cs�Cc&�=�}(��ړEd���D�\�2�Q�|�*���n�LY����v#��ƿ�7-��*�&,ht#B��0���X����*�ɏ�T$��Y��;YF&W�7gͶ-�lV���=� S�f�rn�kĳ�UMf�&.���Lb;Q�{��{��&���&�.)O�r"�eZK"3Gox���|�O�&_�r��G��D#�5�R�����-�?@s�wW�!fU5	�T{7Rw����L3�(�υ͕Q�@)x
w�G��1T�b~¦�{x,^}�u'm(�<���q�篦T �R�����Q����Y�TS��{�a����ȵ8���]*�}a���$0J��*2_����P�H9�ӨA�s(����D&��٬�pk��K���s�1�,�_9�� �}�&��"X�����x��2Y�qd���8R�p�$00��P�*�
��
�_�Ď��vK�#�w��{��Sj�u�����>ȫ~9�����R �C�����5�F�i�Ҝ�`���*����0n���t�h+4^$��#HƏWh�֊�QU�x9�:,,�An���F=]��[��NT�Ik���&�!�_v�U��(���#�)��p���5��P�4���N$���5k�7��X�--y�7UO[���YU�h�B��k�H��י�M�0$�E8�D׍8��q{Ф������������mq�0ի�EaU+/a;��}5)��a�Y����������m���bf���'Ёʑ5Ku$�|�l��z~GUi���0I���%pi���'y�9��`i�][�+��i��}�G�Oi�H0[�!{�*0�Y�q�����"�����e��w|�?#b�d�P_îmRVA9R���۾�[i��B�[�`�������j՗�/�S�	w��kU��z u�l�u4�vQ��*[��Xq�ɂ��~��U:.��j,�7H(VV��"y=��J�Ϯޞ��'�Q�(�F��� Ͽ���D���R��P�v�d$�#�b��Q,��ּq��'	�� �5�Elô!�4�:Ӌ. �F_�ܺԦ�1��M�&��cG��[(��ub�{�ٯ+%��H�'2�I��J����O��M��"7������eR����T8"��N)N���>��6�.g�E����Q�E��L��-O9�����z�A��|�JL]�l#��b�T���{�]_g��ϑ������+�I{�r��KHۣ�
B=��##�	2��Q�, �oT�+�()�n]?J*�������>��?���ݨ�*��+,���	��x��k]�Ün&��e+��5��ƥnIA�gd|�ds�b"�_\ b�&E���e�LAov�������B�N����D=�=t�b�Tf�y�ta�f(� ��}�X`oϞ�$I����M,[*�!.:�؇����[�`rӠ�08��;����cg�%�J/@)ec�0n�˄��JZΖ��E�Ï~��0�?���2ۺ���Of|�t���\a� ���T
��^
�P��m�na)i�,�ɡ�9��&�h"zm=T��>�%�k��vry�QQ]Vx��?�b��gD��¹�p�̸z?:��EF���'Ņ�6HAipe}Y��]QE�Ce��̂҇�E~=�Ca��:�t��+�
pwWVv�&!ȟ]q�+��Ԙ���~B�����^����yЭ��CA�)B�<	���X]�T�GUrI�?V�!���.y�U���w�p���:�;ػ��,���{H���e�1KU�̸�q��r;���H�ŏ
4r�'1�����o����Z�`�*����4w�}Z��M٠2�+��&�<��hGH�;�Zь`��P�Rw��x�l:�^��/���f<1��U]Bk�4ʠE�Oh8?jf��^>��]3���SI*Z��U)�Eq�� sO~���z<�P�4l=�;����$�W�w���C'J�л�}ZoA��m�W����%�����)%�`�R�( A�X�|������yQ&Ҋ���
��ٍ5���f}�E���2�;��W-��m�� O��}���}�HzV��N�Qȱջ)�S�?���!8�*����ldݴT��"M��TL5���mJ;�q�L��y���"@��a="e������yNP��y'g�;|d�?d;�������*թ[-Wb�N�/������{��H��)2��:Ay��67�� ����9�w4�|v��z��>�i�p� ELÞG=���|D����r�k*�����]Q���Fw9����&<O��<��Fx����N0�9�%,���A_~��vYC���]��O�L��&���	S.	�[�����(���mI�%4O��)��=�	�j$��@�7A�����d�>9
�����]��B�X���߹)�ߘ�>�[-�KB�Hv��`�|���R��
x�!ɠ5чf�zC}b=�}����F�P�ǟAR�^��J��M��
��/F0ݚ癧�]zs#@����#ȬC�}�z�.g����T���Ӏ՗�����8�dN+��ʼ(5�Σ�?�1K�1���>&�,�忏�Z��r6�m���-/<P-�'���"ٶ�p{�a�&�Kn�J.�j��	ϗ��>^#�TV�^[�<�$&x������T��`$tッM7��L�35rL�؝�W,ڋGU�A!K�ݪ�'y�����ߵE���pL�BUNx.QK�d���{�!�Uk�N���X�i^fW���'uM�@��Ė�@�}��b��8Nsʣ�)l]��y=���?v%���J&�7��Л�ӳ����T��M�4M�?�-s�*���ґ�$k.Z*�R)�LE]�����Q��*ű�\냐�jl��z>H�͂��tәJ�G�b�:k
�2yp�Ιy1{����:���8��t����UbH��ztg�[��(�כtj����C7���f�bew��➙"�k,�G��\�"x[(����A��M���/���ٞA-)ׅ�BXH�R���g���l��eZmi*,�R{������Bɕ��g����7��և�`�u�lI�\�`�1�˲�#|Z6(u����}f���Њ�8`u�E�8�
ل��
�a@{��Tߠ����--͝O���xn�����RX��IJ=�����Ÿ�Q*�{F�T�5(;O.���ӝ�����n߼0M��oqoq���yuØ,cE��oj�,��p��/I�*�c	,���IR����w��?���A��X��tk�F�ɛ:s��llmQ;�o���!7Wm��R��m��q���xŋc���D���6Rl$��#k����u �7�FͶ'S�&�]��.����o� �Jd�w���SP��p��5d*K�ڔ M�ؿt�t$U^ZE� **��d�ֶ����O��P0aB�����/�>&G�6Nid�� S�I�	��3����\)
cW���TKC[ �>P�t�]}�b1�#�gP|\J!wU.'(RW����;G�y��V��^�I���h �<W�tG�|���uO%�}���gH	�8�Kp��K��lx t�@��()��� ����]cƑ<�2F�jkM'w�ӵ��Zó��K�,U	��M�c��0�e�q������tЫˡ�;}�ˁ��Är�e2�����\�a�ٳ�p&�������}����fY�?>�$�q�.k�����d��dQ�]�שL3,�ҋ�y5�d�tya*�
���T��v��6�[����k��	-�"�=�o9lÍ�iVt/�"&�L��<"�pݹ���O�p��
�LBn��5��^��U�5"�ơ=��jf�r��s>���@q68�VJ������?��ϒ��b��z�3��)q�֥�ˆ�:�w�)Cct2��ZZG���|"z>Jr�/�1a�Gޣ�T�����˺��A�AZR�-V���]��*w`jH�����:��Vf���5����0E�zz:�a���[�+h��0�ݰ��3�
����J��=~�g7ꕪ���&�ќ�����r2�8Yq�.��p�Bk��t�P���Κ�s����N�#�gN�%/yα$�g��lz33����x��R
�̔2���b�O�/8e°ˬ����9^T��5���ģP*��w�I��o⋱�8�z�i�:���._�`�u�D�j��-��B'��r�׉�r�Ɋ��P�R�{�*ӟ���PjO��-�uV�����������Xqj!��d�{�S��&Sև��ظ��^i2��Z��ڌ�?����m��Fy���@��H��97���`�����������2s�����I����y^����$��[��l��&V�_�����^�_����ep.�[_�9g�9��Pr̢@2(�ebDr�ո��Wc���Z�4Hi�N-s�Op��4�X�͂��Cr�MZ��=��'�]~h�%~������"��Y���ӟu���Q�
�,_�`N�v�������[�~Qw����T���f\��g�g��e��;ڍt�@x5�_�iy�B���g���7f��-f��i��ӧ?�:��f5��~�V%R��0$Ug�f��X�����6��'�`��AZ�w������" b���,�#�F�L�,8��Bq��PR8w�2ԉo)U)�`��N�i��+���X_�N���È") ?R#O�dΨ۱k?%lr9tB�#.�4��V��͒������;Ap��/�}?� �N�'������u4��ࠩ�L�>Y2��E0�3Y�d4±�'<�@iT�A�v��v��B'�.�1v+��O��}�i�t�-iT0�d�f3�x��9"M)��c+�fP���x��^*D��G��5�p4/�*��lFr+�v��T�͛���#H�6�T���2���)��R�3uj���� X�lh����]�ߌ���%�j��7�+�89��~����������p�b�����	v�
at��*/K �l9t�_��<"�k�l�nJ>���I��+�e3�T�q�q�A�^����BW[j4ذ�[���6^.�u��$M�g7:�l�s��X��Z'ut�k"���o쒰���� =z�	��Ҿ�C�
\�$��G�pf�6Q�d���.�V	����y=�!&�/��e�#���~y�5S	��2�MT�.����O��K�u6��w���M�8��:�����QwW]�d�a�I�ǫ99Ց�#;������ ������ޖ�)lp�E��nI��e�__��
��^y�F{2n�3�X03K��f�wc$�@������˅�d������װĢ����'�;�2�[�և���GC�#�t*8<�%g�����]Z<i��բvH�*.r�/I� �X�����9,?Xe�"�׌a�/U��Ls	=Ϩ�~;��#v��%̶�K��s��W�����\k;���=���}[�R�b]u�H"�%�d}Plj\�pE�r���V%F����@=y��U`�J8ui�-�ɛ�U���"%�+���M�cCxI�%�e!�e ���A���!%;p�H��f����DDb��ik�͗��e�%�6�{q��x�1W�#��-Ah�f�����%tgx��j��G���d��c��t�!���
�3�"
�@!/S��%�᥵4�1Ɛ|Ã�
/��攛��kd�:U/����o t�R�:^���8#*�񪁃���c{��䣠��e�f�3,�����2 ��
<�;7-|���j�o���wv�d�R��x�r����)�)���� d�>�x�������|�b '�t%3&rZ�̵���,���&������z�
���l�'�nR�2rO%Q'��Q{וM�/o�� �=^Q۸7s_��S�x{ȇ�g�~%B,��ɢ�!8SPĭ!���f$Su/#Q�T���W����P�p���T�)a�z�H*��e��J��hF�A��_���H9�}g����ׇ�j?~��Q��T��%��7rMB�%���NX�����f��Yd[.#����.��iW��˒l��u��ϋ��b��dHDԝ��
g�5���"D /����!=�{81�K�k�?e���݁�Mp^���S'���n���S|���j����J���h���Ms��y�h��]����䉦(v��:�//XJ�����2�=�����(K�0���oR�6�E
��(�vG�r�����u��p��zi��ތp�;d+��\Sr&m�L����zpp��Gjh�QÍ�ŭ�o\X]����>��`���t���S�V�y�.D8c��E>Ś�a�q 	�AD���jaF��F}��2k�0�?9�uC�B��k�w]L�%s1�E���u������;�Ȋ^��Q̉0�u�TwȮo^N�觻�4tw��z�P�%����9IX�w�c1�WrJ@?�]�V��G�Zl:L���<�u��XA(�)��a�A���,��*�+]u��J���W�YX���!��|B*
W�<�n�]c�����3�r!zD���:�|\�G��|�EȞSc��s�ߙ�ƦBl�ԷJc��>���_T���sxc�d�%��mz������+x�\�>
1ņ��I$E��ΠbR���M�L�P��k'#��j� �<�d�_r�������@�&˛*�˒GLb�e��e��ԍ��=�0�hm�r��w{,�j�*4�7j��TԳ����r�{7B���G&3*��T,��u�㋚��Oa�1��y]{�u�~���>GXD����S���G���u�B�/�3"�xDd4t�4��S�s�-�2@n���v��ƒS8P�WP��1%�sU�
7}��I�"��̅�s������|�ho������u�0�Ma&9M�[���pr� 5\��¬W�p{��&Z/���cSؓ���Yʋ��8�*��sA,'��1�zR�	%��X��M$���ŝ-�-ܢ�gf*j�#-�ݎ�f�w `�ђ=�\��0����tc���J&һV�={�69[F"�����P�f��)}0+ T��;F�ݳ���YK������n�3E�9�,�����N�;������w6�O4Z� T���B`����L���6bꂌ�P�^˶��rDX�0o+E=� /P����7Ѭ�^��]���(��GQ�xm���Fdq�*��7��0���7�S�:آ_W�	� 5���q��u�J� �3�P��n8�I�Qɽp&��fOGWD���/'Õ(�>9a�
��|���@���Ei�R�5��}T�a��AP�q��<Nj��iZ6-�'i��-��c_p��w�E]�V�Ob	&\��Ȏ�)�g�?x:��AG�P�2-s�\�Cx���/g�p��!q.�N|�\JԐ����|��Y�_,��}	�������Ƀ�Ƭ�&<�\tF�y�����U0(��G (���?)��}�D�%�/}��=]����I�Hz��(�ƌ]]��zF���(�ed:�P1,�E{����I��b�-@6W���z �f�Ƌ�]��h��bX9;��[v{
*`a g�E�I���)�.L��x�M{/�[A �V����7�ب�1�.�����UZB��"��e�i^�X���������:]a<W'		��\�΢*��6�yb"���]�J��b���+$��v`:'/@��7� �b�7찱��=Sj����Ѻ��O��hˌ��8���z�s�n�daC�X����V�M� ����R�B�s]��	���X'B	�i쉘�����{ń1�H��6xAq�"�	pA8 �j��  AryJ���[����e3R�6�����.0=� d��	�!�I��Ӱz��D���_�;���h^��8ۗ�b���H,�ɢY��!�����rʥ�ӆ���<'A��W�|;�ƒ)�!�YG�K�~%[J�	���a�|���!(N
8q��?pY�x�U�x�0`�~�c�؊
O\I�����X�V�q<���W��H��
T�P���~B�f�F3��u�V����m��򍡜�KoU�'X����3����y��Lit(/W;���bp�>��ܣ��f|
��T/�#�}x�����9�<��q,�F��&'�p,W��c�lUdu_2�YL�e����B�8���)i@���1$O�V�W�DzUS��S�>_�%gn�mb��X�Ee��1C�é/}��)�!�.DTv�}dּ�͝ѓ�@�h8�hE4���ȇ�(YQ$+\j/����6qIx8�_�;[�I�c���mF'�9w���X�G�ǎ	�Nw�����N����p�,ni��=y��PZ�o��"���z� ����W� Ɣv߂�V�7�<���*a��`���'�i�<Nc�����̝�u��xL���#{��!B؝�N����@��M��H�l2
'�����YX�<�*}�h��nK;������\׭��X�	��U��Fg��B����Ç�=����Bk�.bfv�����s���pUy.����W߿����@��e--�����|�l�]�a�V����T"��: ���vQf~�������$�C���h#�Ko�������H�Q?n�����}(j�HƸ�4�n�8����{�LX�"��Y�E�Rآ�v����A�»�Ò'&!��I�vD*�ek�eI��WPk�1__@�`o�%��+��f8�w/�UM*���ݯyWT_���9�Nt�v[ݟ�� I=s>c�������;�𨍦�~Q��r��l!�� ��y�'Ar�:�I�tv�K\���p��)g��ث�B�j˻���{��>>0V��X��m��볅s�섫�*2v\����9`4I�����5�0�'徴X��������j�@� 9��8+.K���^S������A�p���W��C0�����۴�*�43�����Ϊ�������Ys�&Ћe&|'q���{���Y��:���}��7�+_�U�Y2���.�a��IZ�F~�N���^Ԧ�\������${�TB��)>�eY�64���T(ܕ�DEIÖ�Q�f���{x�Y��d,�؜����O�v	 ��Q]�c�M����zZ覗ٺ��(�*�ʼ�눝e�NKk�I����m��'��\"�a+3W��Jh�y���) )m�0@G8��p�4���,dC���������q��AL��,�/�.�Yd/�xϲ7���&�VT'�YY]$녴Z(@>�^*'���uhNƭ�G�2������"4;��E�5S�_[��hQ]��\����l^�E y��F�TV�%s��WT��e�}ozO�<*�	dY�C�2��������c��i�#�ؽ�;"�iN�YOl�!�� &�▌Y^���E�H[�"��2-�4�b�G���}ғD�FuS�2cD�cAP>��)��w��'�GY�i)�fV�o��%��0�i������F��]7h1+�V�H'��I��D�i���I��T~�Y]�d�Q��E= k(�z��C���FU���'�M��[��4Ӊ3N��۸e�Ԧ:��m�֗�l�Zd+�"v��WIֈ i��s�dǆkq
5��
`ҷ������!����$T/e�����p�ǥBBz����PJ�,zE��J�lA׳�
\lݍ�V{s2}a���%�o]6�(4t.����Ê��4���5<�1c����]°X�!k'��lx;$��1+��?<��?#�O�7r�������YX,���U4��A1oȚ�o�d�P��L!$ݗr����� ڸlE�i��H��2��I� aŜ'��m�ߑ��_�]j�2acHc��%��� �=��q����w�J�К\�6l+��0$�w�5b�a�f�K�HX�:��Sv�u|��9�gÓ��K�=4�����j쁜��8����=�_+%�!`����B�qѤ�Л��t�K�b~w����Ɖ���i�$��7�=)M�_�C���۞�,�1�]���a�=<$�78�j�	'!q�OB�����`���zt���5NIǃ�g�NL7`�DV?<�\mY�~S_�ug�3��_�	���2g�^�5�P�;��435K�&�i�$}2b�H�ۡ��!P)I�~�P(��W&�������~�����i\ޥ������5�G	����'��U��CxL�K�6~���+b��`�8��Wy�L�}�
�	�B��s���g�7;E���/�A�u{ڢ�jr�>�����9���j�!nZ����|��N���")��b�Qh	��2�E�1��r�p	��e�/���,B�l����9���
�������� o�O��c.�e�c;b�)g# d��M�a�W���q��:�I�������|��B�Y"9���g*�&�;F�BqC���#��5
փ70�;��/�a����_���\L�̳���Ĵه�xj������,Ŧ��܉Ld5�[���8��-Bi�99^�ߥl|���'C�[WʋU�D(�hGc�S���&��!-!ڍ����h .9!n;Z�L)5����NX�<?dow������Se�]��ㅆM�Po<�3��]gO���$9�ZGW1�1��2	�f�zע��l�f���HE�o��*KT���LRTm���K�G�Sg��v��3�S���N�
�5��w^���J.��R��T;Հ_ ���A0��D�7C$�މG��R����n�zmG��ͳ��
��󥷬J��Z�В�v��<�xy����J�p4uEv���B��+0��6�byӋ&��~���@ds��<��I̫
�A���ķ���� m�^���K�v�	ӏ�>vY2W�tK8�	AA~���kMY*��K0_��;s���-�[t~�G����/�]9S�\ti[=�a�	1��!�j�t1{#q�	�w!�KA��]��a�/�$�A�L�&B���;ţA����Q��I��ӊ�{!�~ %si�?��"B�.�~�E��+�� ��?Ç�/��i�	@�'1�,y�.3�:)��Te?AQ� �?��u�8������Vy�\O��p��Ϲol��p���|��{��R6�KzZ��/�[ ��&{�_ʀ��>Ȕ>��gNK�W+\�	\��e����^0���F�E��`~xs=�!����mk���^�69�,�HzsM�/ޏ��:S�H����D;9�c��īI^#��_��ެz�ʗ��vEea"�E7M�^0=W��BW��J���ϓ�&b7s��/G5xj������l����c3e�/7�q�c�â
&c$v����k��A>L�S ��ú�V�Y���>!ڧ��~G�~�-�D�1�g�Wy��P��Y��n�I��/�1�>��*k�Ǭ3nb�����.}�{h��1]n&����}���Ё)o��
:�g,�� ��T��#Y�6&��  Ld�v*�Y�>���������x�&�k��S��*���i��TA����hf����>�D��<���&�d#�:_1�� e��!���:͕�X�F>=���@��o�����ו@^��V����v�Zw�"p�n:���MLKO(��M,���0U�_bJ�i�%[�d��K��G�r�/����c�N?1��n~Y��p��2<���x}���d��i.����/M�^
�� V�4�&[<O	_V
������-aR!��ꜭJg�p+�Ҥ�ꂃ�s܅@�Q)<V5��u6D/d�q�O{��:ҥ'Ci�n�X��d�E��o
���σC�E&q�R�ʬ)�:�?@n��֯�V�b�~f�D�ڢ�_9�����Zo6�{Dp�0�b�D��@<�[y�;��&����I���Ł��7�����K	Li�y
 oqǛ8���l�c��	w����z
�"X�",��tk{Rd����A�WN����4<*M��)J�K��Z�9<SD�����ݹ�?m��o��]����tP�@R�&&���ˉlC�i.� ��`��`^xK7�'��M�T�.�v:�/w�u�Xh�1 �T�l'������7���a�R1��2� qs�"6yv��1�4���uC��J;N��16�qp"��h��!{A�m7@�F�E�hwl�@_vO
fi@�+a5H3>� ΍��s��he,��	��������-�D��M�r���Fכ��L�rh���E��ԂQ� ��e��k1d�OF�};C��(�`'Ȧ2zL�2�+ֱ���:?'`7� � ��E3C�P>� ���d0&�G�c��ݑ1\:��������@�t���3S�����FH��=���^ڇ/hrr��z3x��j9ғ��7�/?m5F1͚O�B���2:l-l3'S����$�gnޢlc�p���f<.�r���_c;���dĨ~��.�Ƽ�x�ߦ1S��Z<�o,d#)cl�-A԰�qj��߬�I��%��c쀕�*��!�XN��|��h�Ei�m���#ͣ�y���{[@F(=�ԟo[�{h]\i��	������|V8`�I�0�K`۲E�v���T�ec�`��i���(J�����\!��&?�����ד|�K)�����UOZX�~�Ͳs{�oIyqN����Qz%	N���u3�˟ԻO�vc6jh:p�9b��R8_�N�}���B\�Xo��T�Ǫ��zÒ�}Z��i��r��S��h��ip�}����݊�fǁ	�׽Q�p�a�����OUW�M�K����g���3�4����'
B��t�ώx\�vZ�m��3Q10k2-�m/�̯��E'��Z���P��i���]�ғ���G���de��H���hQ���NG2D�gf�JZ�[എ.����hs�O���frIspr��I����3⣢�5��<�OK�nFX�V�Y;�I]o�	.��ե�K9�c�Wk.i�#��rD�����g��s:��:�R��JD����&˼Q�H_E,���3^l?m��$��\o�=X*Mx�z�䈡$��ҨJ8aV�D�B�|��gIN��M#+��#KeV�uh �S񨪝YƐ�&3�D��+,��~ch@�.Q� �9�l�Z�`#��Q� ��kՠ,��=�#�nwjZ�l|H�EO5"s��z�W�6����.�ܬ�P6ާ�^����AcLa�h/��<�}ʟ�m�Ł���K����`V���%��C��xt�|5i*z(g��%.�����i�(q�8��]PCq�v+g,��9��U�涕�O�'n��}� ��7V�kN&�G�e�i�(	�^��k
�$���j��W���s�ta����q���@~��Q۫�5�L��j�~`.���]}���l��oYčP�X���(�'dN�3/M��?q�^�/V����������<j��V�4`Z���;����T����w����`M\��@��S��Y�B�Q)K
��]�߽]PH@�����`ң�*}=JMȋ>�t�>����qLNb_�a��X�0��9g�������$)l>n@��E�0�V �x��L�T��ae`d��v��өx��M9�CTY��޸[���am�f�Lj�S��)b���׉H����6)�ϓ�*��8�Om�)��瀫{����r���=$a�3���2��Kw<Wb�dXhmn-�/�$��@��㬢tK[Zb��<<��~���5*~<I�����߈��-����	��[ն�.[���
V�t�+<e'N8�{�ˎ��#�.�G�9b��+�۝�? �S�:� V<킶R��M�����դ��]m�,,�E܃_��歕�b��;�
k��R����w�p�Z���J���I��
O��wQ�o��(S8$eEٞ�����pn�yoW�}�G%�r�!z�q��|�� +:EJW�QJ�yJ����T�K�f ��J�R�>�ı���i[-e��ћ7���L�dn������}on���oć����J_v|2)�����c-�0Q�R2���Ƨ_�{)�b���J��:̡5�8V"��@G4.m�w0F,O�po�k7`t���֬�9f5~���a"���W��xw��O����3ED��M�R��^����1(T@�y�%JT'"��Yt�M�U�D�1{>b�|�Ώ��`�C%H�j�,����vY2!]�\��������6՗��h�\�S[(ք�Ƨ��U#�)�C�yԣt<��5��3笥V��W�5�	%�Cn-��GY%*1K��˂Q'�Q�s�4I%;-�����4P�]���M�)��aق#%�Q1h&@����a�����t��/�Vx�jWm�7"�8�C�ʅj
y���*�}ir]�/{%�(t�k�a�՞�u%7�݃F���?bSyǣ�  [����xa($�U7�
j0�J��{��}B���X6@�B�� �Բ�Q�����^�\�ߌ�=MAp3��k��) �Ѝ�8o˹�Mcd�IAD4i�m�׶����o����#���Ƃ���@|��B��c:�R�zٻ���p'��"�k�Qw�����(N���ivuD�&<�1�vo_C�S6�M?��-�E������|�DZ��i:�!�AHߪm���E�lʌ�L�kW��z��� |��P�P��P�e',�I��R�W�]��hƿ�qMd
�&�ն���m���F�����:�����gƙ�n��/����N���ח<:�����D��`��\\!#��byH�XD�ߠg^����kv9�N
2m��׀z`�C��΀���L��Jb�}��Nq!w�'ًu �Q���J�f	�6jw4��f��=c���`���o3����j>]���p�5ؘ�_;*2�T�]�P�+�����r����Q�||$��%�M��S�p�@����Mc��� G�ϝFE����Z�lը��g?��C��y_������:��'fǻO�S��\0�DM�X���ĕ���\_B�
+��+�G��P@�˵�V�sb��Y�ݽ�	��gapQX]��dYJqgEL�X�S�qI����_��e�����1;�t�d����O���	q����	5QY�D�AT�
�S.��R�F����o��u���PM�ҟĨ��W%��L�B
'�/���0�0l��s��`s���ך�c� �4R��>�Tx��ƞ��hNo�*It����������e�b�Q*�d,ѻ��瓽��i�,��@��0�Xe~m��׆h��C'�k#>�hY�s�8[i�^��~�"v�Q���g_90����2���H��O�oN�d�R2��N�O��������!�E��B(Ph���H�-�n7Ͱ3����e�P���<�&a$�����UfrtK���k�Q�O�8�zJ��e���}g�����]ώ�Nv�Փ(�7x�v#�q�O��תN�HS��"]e/E�
���RY�F�6/�M��[7�F�|����iI����s-Mѡ����0���_y�Q��@��������̄h	3�q�%*S����_�5��\;�����O��~x鞶-�����գ1P���K㶛����ȗ�Sz�F`������n�䶊��v8��vxڰ�
	�/�,6���\�ar�� ����h鵐�H��Q���⠒��E��y�P���ճ�(7�k� K�D<߲�r��ҹE��j����JNj���ć�\K(П�<>5V:lU�[�굷;�� D�ʶ��l5�����`� YhK�Y�C�.z.2sq�1��|�e�|�2>^�p���n�F��V�ت�џ;�9L��ㇱjG`��`��Av/,��v�F�l��~�I1�&�DnNqD����a��<���@�=��$�7��k������H��
mF�vy'OK�T5��ՄJOE�_�U
�M~8ٟ1y�zAo�,�QEG�b�~,�6�R�ӊґ��]҇V#� �.>���lֻB�S�����& �6B��q"�V�zhCѿrK$N{�z4n��j"��	�2�1�1�@*k�
���Ck^0nD֣����qF�����Np�t� W�p$F�k��Y:�|����/�0�s/�u�@꙼љLm/��=�b}���rd�<��9w��-�Y�qS���d��e�W]�"X��"�y\�8*�~θ ��9��%��U8%�MQ�N��{�x�#� s��m�Wu�.��)z��4�գd������$��c2*�q#ĩ�#Y���:��,s ���f�?�נpfc��N�j�7�Q9�C��	>zB=�H�J��|�� Ҳ���N�I��`$xV��Bp��x`%������~��6*�v��|��Ja�]$Z^���\"��gN�6���L�n�K�΍�=��� &�X��h�{3�#�1#W��'Ov��J�[�x��Q��R֧��xx��=o9����7����>9XU�jT�~�G�(X�1�\m�����6Ot��*�4d�m4$M!��+��TF�ϓ�D��q���#�4��ek��CC��#fq�ނ%so�ǱQ t0­�Ej��9k�'JF�&M1�y��#n������d�PKu z|�Ʒ��uh
����V56�C94��lC)�Z=�|t�7Z[Q��W�S��r�i2�P��_���fJ���e-�Qk�ƛ4^0�Ȁ�=Zژn�[J��*����M���V.�Ń�!!3;���D�x�7�0����)rCz7�{HP��<��uX!;�)j�r۶����⥓Xz$�Ww���^��N��J����lZ8PGk�|��������Zv���P�F�.;�3�̳z2��I5f�g��U�՝���O*�9��֗z+��
�)�n9d�]��~�[�덥n=�02��K;����9��y�A'���+S=�'ݠ��������B-��l�r�㻖�*T�<p�yKX�sQM4��=GO�p�zӻ��S?5и�M���D�vQ���u�F�9���w�MB��fl�+��E�O̝�6LP��ݣ[r�m��)z�S�q$}�R��RΑ�4�@�sV�Ew��I.��M���)�KW%j}�yq�4wn�ٸjS�6g��tT�}��V3(�2��s��T�� �̨{&(�:��Ԡ	��t`ߟ�B���+ԂT�b�w�5�)�W��*9�­���f��U����R�%qSz`sd����3�u!�.R��+�v�����bD1�n5����TRΌ߉��s�2jH׌~&1��wf�TM-�P���ІFJ�W=V���̓�$�9#����"/9�)`�u��������S�/{��.J��r6��g錻� l�3�<��_�'��q�������z���:ݼBV9մ/,;|���m���Ln�R��w�KtH��F[[�VAs�M3j�>��k�Qπ^rl5���Da�hT���%���&)�ڵB�
��	��PpVv�:O�/eL]OC�L��FEJ��u� |gp[�w�o�(�m2� qck�|b�lD��g� R�����],�9��z�Y Bܝ[f�2W�ڤ�Y�K?�t���6v�7
EyK'��-���T	^
Q?k(H�}��}R�4W����Nлo��1E�IV�H���|��X���o�aѕ(�i^�=Y�S�ZoG��D�o3�"OM����^�E����x��*b�)���2
�\�άƙm6$�jUCx���O2X�Ϝ.䢂�Ӽp��T_��`�o�_
^��L�A���0�+q�}`:˾�����O' O��O��K;�l���_Z����m3�9�d�h�s��V,9��,��*~`;�-�K�a��B�T�¯R�5������6N�IL�*@B�&��҆�o'W��*nz�
��
�[����/�B��R��J�G���w'�CO�=�x#`�]�	@rT�ΛHT>�Ho#N:��h�6����1i#3��w~|��tpjP���Ҍ,`��&3G�W��>�{I�g�l��ކi� �𖢲|��m��_�Ί�<,�t�x���^�3ꋬ�~�[�j�{��?�,H���n �$A�vI��E�ſ3v��w�һq�h0�p�X�@ �ԟ*���o��9{��x��>&V���oɏ3
ʯ��H[	���-#��g{�� �/���L[_O��/#7��Z��"�h_gX���E������s�iOzK�,�yuP.�~^����C��Io���%[�	^�ҙ��[�n�5߽����t���{E���1��~��5ߍN���o�l�G��Dv�\_��
��{�|�H6�pF�	_�_W7����N���*�����*v$����
�˙�����i')|����y��^lv�]��H���H�`��n��`�Z�h�҈_iUY���hg��=��|�ck%l���ש9��t�F&DK�X��7=�ٜ}��P�r]����hZ󁄣�{b���A�C��:2�m��Yq"w��c��ybS7�u�E �l�FB&|���}�t4�?���	��[$ � -�.Ѹ<w��߆�o	�nps��n~VS��(���Gs���������vG�����&C��;�j������m��h�u���#)$^��|c�������X��[d�??���<Y\�ɕnͭ	+C��t>�n��c�k�p���/(W1Hm�i2����|��x�Z�dt���Q�r�;k
�����m|��,�!SL���4��"��4ű��\��L[��m6�0?<?�����, Β�fl�ĭ�&��"�1m�
�¤�sj n�q�V5�qa{t2t�G�aM�u��m��)�mf/���CT� �㙳���P6n�ľ�%�9����Yn��bځ�m3ᷲ�K֓�~���]�Ű_��>�#]���,8\�~?Q�0�G���u�E�E��+���Q$���0.+���8��q��x_�+��d&�e_P���ʼi��N���zz�*�3YU[.�o�� �#�r��C-��3�"O��$�l��Y�S
杗�՞G���)�*j��5�T��=��Dn��e�l�Ͽ��8��mKK)E�J"?�����a7�������'-+֚i� (-]�b�h�p+�|h1�z��WTSPL���p�v9(�ѭ̒jݬ��JjYi1�Q/^�q@��5N��x�F}����p�5�፤�a���ĐG��|xAn���������Ff�i�׳��g�Hyg\��ԛZŝl��'�p�,|eo��1Y�@nrl$��X�� ��%��1�|~wX���C�*��Y�}�<)O�C��o���EqL�=�L��W/?��aL�{�{!{ �GU�}6��m�����M�(1�B�;Y������-m���bX���%�K��%��O�.[u�Mr{��� �R�k	mo4�:�`}�M�S�����.ѰI�K�H:�\f!�T�Gs0�|���b+��hZ��A�`�R'E��6�n������enb�5R�8|R�������?28I�k�����)g �ۣ ���6�O/q=mo1���{� ��h#����a����qܷ2�J�g0�gs���@F��ި̽a���j�L��~�p�"��)�]���TL�+����t'����9<eK���iN�Tg�-�Q9�h�w����=a �y�����ˁ�->�z�"�˿��2Al�冝<k0��p��_fpa؋���ӊD�^}Z�˞ff}`2�v�k���y�R[�_S�Ѹ�k��φ*�Qu�io�f�7{�d���-!�=��i��U��j��TK=�6��Cj���
���L"�0��'�N���û�E�_�;��g��>��a��eqS�h�u�麆
۪I7(���^���{���p9�8�mR�pe��Y���A��iC�꨽UΣ18�-c�����3l2%A�=��a��0cz'��T��b����V{��lB��5����!q�ixU��,D�l5�=|^����������%�1z�-���RCE�u��b�7y6�
��{�C�/'%�O�	��Ϯ��!��>����m�>"*���^����.����gY�u{��x>|h^���N���8þrC���;/�����Glӧ�%��� ~�h
OWK�[��M��8��*7J��X.Z�ؠ\��P��
an�:�z�V��L�54N��f��&Xƍe��&��\��bP�
<���Q������1V�9z��p��2��m/0�uwM�(^���m7#ݚ�j����\ff�~��VFA��}�@��]7 D}GI-kd~�+�!=��Q�ɖ�Ζw
�E�
��v��q�7�)���X�|яu�����^^���,�\x�(�R-~;X�ʉ�x�FZ���
&��K�n^}¡n�)��S�M��;�����̾���j�q1
|����6��b�����O	��a!zk�M�~��{�#R1�N�$�l��w�0w�{\|��kboD�v��y��bL馇,�+������@�����.BVWZp��9a�8�cĆ�J���h}�K\bq�u��c�&��U�O�@,�1�SG���9�<��q�)��6�1p5
J<N��HG�9Æ� 8��ѐy{��-�L�����]K���X�&
U�o�[��<�@
d�	T�xנ��Y"$"x2�-�b�X�V���9��$<��!q�����.螽F$����Uy`]�k�C(��j��+�YEp��%�4�&,џ��<EB��ڌ쾯�2�.\��Z��mޗ'��U�M��#�&�b;f�T�0z�SyX����ŧ	�T�#C�ރ l�����
=��$�M�i/�L�M���z�gmy1�� �.35X�K�2Cٝ	7�₇X�/i.;� ���M2��Y9��(|�;|R`�ԕl`5�C�Q�j�E�GP�m �m��[L}�ȱ�>J��!BrR��ޥꌦ`�
1tMePL@,�:AM��S@
�r,>�;W0tyMt�N=����9�$y���K���[<X�|�'��kK�/��O��c�	�B[ׄ�P0Rt���C�Q� �'\[�h�]Yn���~�ϛ��Ӎ�E�A�āA���2�Q#ȱr�r������3\��{T����*T3{�'���Ó?c�D#+�v�O�^�����xL��������zW?��j�lv��eB�k��@����CZ�x� �y�	��L���y���jO��a����7.o��K%���Tà�C���ȵWq�s%�l��pΦ@�y�4� ^�` zE�4R����_�������ƺ3�|s��F��T�O/��}��H�|�~��=q�?�Щ�������^jY��X�+�)���3��l��^��>p:J_z4ט��z�w_4m�!��t}�Ռ�{U���׊�C _O�nsF�ܢ�j��F6���2��ml�=r�qE�InZ> �����������/�v�P�+FYm{�_��q����H�$�����J����/M�E�ŭ˞]y4u�GCDpsBF��Yf��${�E����s�1	�k֏�����v�f6Z���[�(�.c-������|��s4(^-�@� i��xわfB;�<h��E�]���fiDv�4�t�����W^��H)Z&	6(��1T��Lm�Bs@�KQ �Vq�WP���1M�A��6�C��#��;���P�c���UF^�R�p���z����1XM �e�@������C����a���}��'�+�PT�ѥ�9M�?��h��n���/�hH=�[���Ft0�\�������������%<�q��T?����Ks���Lv*zB�)~�]��dr�j����-r��{ΥYM�(������}�D|��5 {��W�;(iUv]��uE@�?u��*#��ϴ"��gKT���a驢�X�x'I��5>=��6}��GP�
a�nR�n�%CP�z���^�����$��G�c��ڻ�;`N�4���;NL�j��/��F�O�d�]�`y�F���%$o��(�YA��#��V�y���ئ�=)h; 3H_��k�r�Q3Q��%�����$}0�7���["�S��@��Z��w~P�K��D8M�UX{E���dQE�f�i�����Sw�Kb-{��h���a7�2��B�C��'���˩�W�lFܼLq���B�p��I'k�?���Q�{�o���a1rbE�(A����P(��r�qR�̽^DsL���G��#���L�~��r�J́2V6~�@��r�h:��b�W.�OEl��',.*�NO�<);���%u���?�'I�{�Y������^��f�o/KuNOJoi�p��o�Ò�܄$�AbO$�9����*�d����ڙ�D� �����P�Ѱ��%��$J	����|� V�I���;Ynp\��V���չlE��t"�m���S���	tŌ�`��M�v��2ξ ;R��a}���+:W�Эx��Qca�AñV��֍����tR�Π-�������`V����3�ny5ك W��Y��m�-���K��լ:ȴ��}�̈| ��~��z�e�dG�����3������KK���fԥXj+��T����J!͞O�(�a�lJO����1ݹL�{������`���Ǆ8�	gG��fЛ#E��*]67�R� ��_X�	�5�I���2^U?4O_9��V��a�U���/��Jϫx�B*rB�%Հ0l�^���\"����W��D�q��y�3A�
��ʧ�ֵ�:�9�)pPeSB��z*��E�G6�њ:t��dy��/�Ee��DU-�n����M�����$��i%��(�E�)�r?���6��RB��ī�X�}���o�=��q3񨓣���3r�}5�r�L��!�+��WG=e�Q+��i��zx����	�Ӌݮ�1U�Fwݏ��fC��"�k��|��_��e"e�r'E��UcĹ>`/���62h����Gl����ŦÓY�}إ�AG�#�n���I��� �<��_�A����(��I6�J�{}\D��L�Le9lAVI*��<��1�R�O����ݼ���J:�N�=�/�mk��`*E�<R����Bp}tFN��'�cmo��^T�Â��������{��0�'6��Q�>8_�͒�O��݁�k�'HПns%^�r��+�2~��l+Sá'��Y��-��ӏ��,;gͧ�d����<Et�� L9� ��V�Ő=���cD��Ks� �'����Y��|�D7��
����JJE��C�;t�q+y�s�
��Uw�wx_i�먮S���ds��w",:�׀�a��0O�$4�IA	�">�],��������*/�SC�=��I�am���QD���0e�O��\�I���x��|���2��D��f��:Qğ{�D��E� �~�?5A�L࿔1@�rs��	�D�c�^ضd F�����]���b��!<�w�E⃒���3f�#�N+�Oπ�%���s��C��^�,��k��9S�.?>��5*�qu4�~�Q��5��1*�vn:����KK��� �wH�kn�nw<^j�	�(J��裈��+��?w��ƙ�v�d��>���(e�Rw&s�f����t�ٵ�[O�p��.��T���j�\����9�U"���Ort	�p���.��i�l"��Xr���� ���A#͑\5����r��7=ɫ�2��Z�Z�jt\i3i9\�P]�*/�9e��P���(���aC�����1`�����v�xi	�Rѹ�@����x�ʄ�j:5̡?�O���a`�8��b�PIg֬OSĬ��	�b���.�H1��s�v5�����8�.O����U^e�+o��:����g�p�#,�v�!�A����lΘ�vܱ�F4ַ����V����Cpv�����.��=ԣL�*J���mp?aǮ&)�Z9%E�PQ��"毉]���!�M�G�"��H�� ���-��6UJ=����Q������v����k�>�&�s�V���`��_�,��W����H�s��%�]��}�0f9z�S��y{�Mt-Ĵ�	����Mz�Ȅ�_++���\	B�Ԝ� ���b�cZ����$8���/zg�sY��r���R	��RR���i����)D�o� �1��뽠�*�9?b	!RA�_u�!�aOBeذ�ɏ� F+-@����(�a뮙Wv�\G�{�\���?��P"S�M�͗8��~��a�YZ�+N�!�#����F
�*��s"J��6����՘N����0���K�p%�}M=�vw�t����Ai����������e�5{��T|�4�۰m�T���o�Ƌf����\��,-�9���m}WH��7rg20WR���0c"K����l�7�D�t�Ǚ����m�HG�w�WJ��C/u.�+��bl�����6�d�Nmw�� ȓB�6��H�����\j��>m-b�{��Z�'ts!(� 0mr~<r �MVj�P��LOP����"�ײ�vՎN������e��s�.c�o��ɰlo�M3Y��rV�@�h�.��)�_����n�!���&*����wЌý�H�:�Nݟ��ġ��ߜ����C��6V��pm�KU�U2����]c�y��l�J�"s�R�9LI�֟��EG�/�.V
��f�+�ˡ��$��?aҋx���SI�h�	��yiR�ӮB�>���]ճ�wzk��7H֤�;;	�Gڿ��QA�L�u� ��AtAkѤv��w%��Sӵ�Q�`�U����FPm�n�^�ti�$�j珶NE�u���3C�~e�o
.���C:�Hީ��E�^�Xi��gx�����G�T^+3'3�v��Nc�i��z��^g�q�1ˍ��Q��X̐��;X2�����*A�"�VQ}&�{��UT9%=�!r5�~Hm��1��1tw~ވaK����t0�"iw���@���2@��d/�9h�!C�����b��_��HP�ZO_7�3�.����<����V�%I�u��6�ͺ������M�3�ʇ� �<a*���	,��Tܬ~ѯ<�/�5ĝ�����]��߰C(�1/f�I1yK�Ϻ��|��.���I��'��.��<
5]O:_c\7����}!B|Wu������3
U�9Լ�a0��J�53vU{�!i&�>S�L"��#�iJ9r��E(�5��uGby7aܾ��6�)�,���d<g��@�1B��Ct�{_�3U_�m�m�c�k�~|ۍ/QI��ڕ#�s�<����m �����ݦ&hS3�W�ε�-<$�t-�e�`����Y�o3߁hQ��y�F�_���g���?���撐t��i��E��R��O��\5���"ӷn�O{>�`�%P�*'���o����ҕ6Gaݟ�0�5,m��>�3�B��6�Y���j=G��}���"y8���0�����97Jv:Yl>0�/�ˢ\�6�r��G��ߠ�5s[OXuZ2�	�,a�QJ���~7�`�>�_�<ײ�w�o))�ω�`{�K�>�0��D�nW����BR�EJ�nJ��w���RQ�w挽�Xa.:"�}�(�T!�K�2#ڼ(FAewI���ٯ��ҕK v�WTU"8_��X�O���ӄ���$���P "3k��ʗ����]��KF9p߭ �WÛ�G	褓%a�����i������0���+�B�7cl1����7����C����?O GE���	<�L�c/#}���u�;�ncj���+�f2t�L�}"[;q�=��VD��M�펧��Be��T�qY�S��3_����5���C�ږ+π9�ET�K��:E���/9IK��T��&�2Q�4��>�ț0V�ww����i�&���KX�Dm�ʩ[
�P���>�����K��N�*�Y������6i�?d�t	g��p�g��E�P�c2!�Y���Lh%�^dŃ���m��K���~@&�'�>P��q���D#���<?���F�����89^��T2
��v�QǨr\�y�}f��nN�E�&0�����؝�jl�c�d��?�"!`��\��WI<����g{��eO��Q�7�ƀ8I��#�Uk��`z���hu^#���[k�K��ղ��W�p�������y~��Q�{�y�9�#������V{�-�:G��np�5��{S�f
8�,q��ae��)QڅS!���sA4��۪+�}z��s�������f�e��j�>��o��F��>À�t������p���T�Fu؜t�JD���˔N��O_�{F���	��x�� )���OƳ.�.���7��\b��C��L,� �a ���?�\�;�h?�Y��E�:���@����f�)��i��c��u�zܢ:$���&_a^Р��P��*�B���Z*|l�<�z���)Wޭ���=;Cw��<��~�L�9C�< �yI?G��</.��_X���d86�4Y��1rΪ�b���Y%�g�:����B���^pc%\�������q���rm� }b� �s{:	��Ҏ��w���,�b\��HPak7��������K�#������V��z	/Ū0M�o@��;�=�����y���[�=��	@����O�U�R���c���0\]����_T��9���Lc�n�8,g+��w�b{zV�M�5BJF�'�1�I(��1�_@R���)�br:�ʊI~$d�Dc�=Z���$�|uiO�c���A��)Հ�Z+��7���ZkM���ȉ��d��һ:1�����<���o�Zk>�x�3��g_�b�^�I)��J�ƹ^)��\U����7�]��J�c���� 3��Ʉ2�:mfrj�)ÔJ���%�*<��f�E�r-���܊�粇֯uku�yj��I?"<3vܸµ�D*�����m�:��s�
b-QP�=�E>y�&$��f��+����Q����Æw��y�d[h�~L��^�;H�4g
d ����9��{���c��M�d�D�L !���)�s'\�S� o��g��ȍP�4?>m+���0lf�f����#h�炿�¡�O�Ak��/R�'OH��0�M�Lk7-��m/H����ߪ��9	�[��<���g��;��&�L�0��P�Vp�#4ǎD��#�*{|�F��	�2�S��)!��'Y�Ǡ�����d$F�@럇1J������ϫ������<"�W~hS������T�_�����i�Oa��v�IQ3��-a���vD���- ������V�?4�"2*t�!�u�� {����O��K�ѩް��9bT*Y[�	�SR���ƺ���U�����[�O��Y -$�P<s���(�>���m� ��w�|9݌���,�Z��O���b]�����-���<D��Pq`#���n��K�TO��� [N8V�l�:0g��A�=9�99�F[�^���bl�[��jP�o?3ZX��k��v�m:O���&I-`b� 4��%,57��� �u���nq�O�#�RH�j])D$!@s�Z�8�PD�#���Ϗ'7�C<W���]����Z#f�Zv,S;[�kMb�ݵ	�"6m�R�@�X�N �bHl'5Y���������/rb����gn~��������kNz�4K�1��r�ۻ�:uq�ɠ*~�j+	�b��e_x�N� }�#�".��?�R�:��6΄_��fX�d��zJ5��ţ7��C�'�/㳌�^F�qfPGVțȨE�HR�s�R?���B��E��Ώb�:���=�И]#`}���3�"q25��䘳Izl��G6"��%5F����o\�#����%��k����i)1_�>��j U+��0T�3~6+HV�v�L�`D�7ncU:��틿|��>�2dGS!_�Sg ��s31p�Ў��a���Q��b�X���];9�j���1��Wt0O����mʔJm��ս]�� >���8T�6W�J��hd9�B�(l�P~�[��E�@�X��f�
�MAF�Bk+@��r��=J�h�����iqe�ۜ{�2+%�hb�1̡��5DDC3\����-7���?���G��%2��0�HSiRy�ݱ�a�
E��e�Oʧ��]g�r�:�'-��/.�`F~="�wJފ#�m0C�XؤMl������6$�g?kw
e����q[`��ioW��w:�T*�Wy��Y8:aC*�\�Ax����22kPaz�*�))i+�P�^�Ȫ�]iS.���'tG����N�2�#�C��q+��@�*�y�T�����q�>���qok#���)���?��ɛ/,;�&�%4�u��*z�T�0��O&�Ǉ�Po���O�c�G��@��Tg�~��o#�3��W�����H���D1�Dw��0ǿq[*��Se<\����� r|��ĩm$��R�Q/��b��)/�h�3**z�%1v5F�"�J�	����䩆���Z�̓����Mh�'���>y����H�e��z�����D��{WVor�Ff~T�ڕ�m�8�B�cZԤ����dU&�'�fCB�@("�ʱ4\�ȣX�ѷwhފ�2f��_ �N3�[[]�خH��W��^�`���d}�:�X�8�Ț����}*'��FƟ�;!�Z�s+���+�m����V��t H��8M�<���E��d���t�J�Jp��b�BQ���KD�NA�DŇZż1�:��7�lD�S���?&��~�pf2��t�|H�g?�)cV|`��F��]�46�i���E;#浑ah�1����J��6L��/jXA"pη;�O8�Fy��D��1�@�JWvb�PℴYzO'�B;���#Ћcc�c=���7�DS��zL���ŀ ����r�t풽50��6��[�?�iU�l���b`.��iD]�>x�l�0%�{|��Vop U/7sʌ�W�2��2z�\8�-���B�	��U���)V-�%��XT�|�[�<��Lg��*i,G�m��"7qP�1�?����m:���%���L�r�{s���~M���KN�r��{Hg����bl���� 7�|��(�eR���|�~;��6ޚu��>!�؞�i����Od`�W�-����'\�����b�d*�ylj�}k��k��E|�HF4b	�y�/�X��3*����]G�cM�+e>]�6��zE`�H �[��wKI��a���h`)b��d���|�]��$�� vr�`P�eb˨N�b�f���0��-���L�W'�k��.��9���Z���I� ��U�����V�\�2��q :�'�����gbZk��j��j��@q���#^�?����Oً�����@m��ij:}7tT�I�1ߔ� �y�H�7;��R������x�5r��\����i\s�c�Q���|j�|fY{�9z�J&k9hē{���L�A��iPF���U�,��eW�Eѣ����?�D&�'�0�
d�h�7�1�meH��	���yn&��	*��P]|�0{X��.K�\/8RY�%���􋮄7NɁ�-�#8_���>�>:V_(�LXDS��J��w�
�=�5�X�0F6�eA-�r�v?!:��b��k��8ڿx��A�qyd���QԺ��k�e��8���E��)ݭ�]��*�Q�EĖ��I�m�s�EfC��H�^�iFKDƢ#��ގ��ӓ?��Ul0�6��SΈE�(� Z��CmKJ�<�/B�X6��9���> ��g),3�-S�ǀ�C�H԰٭�b�\H��k�� �̥�����������[�KDVxZ@�s;XP�S�`�;�@HQS��[R�q���N�����{����TU)�\?�-y���������z�R�&�!���,�+��?jh�;��b^�.�����h��s<�Jӛ:sX�^����3� $�6�Jl,KE%���'��%9Jf w��]w��U(���§�e�FF����[{4��ٰ�)��">���u��uٓ��wu�Ћ&y��djؐ�C������w��D���ɕ�J��`yX������(�/{C`��@&������x<m�I4"JA��D�"Ui��<�Q~�����5w�GV��J��WV<SG#����
�4�>�:3y���`K�؋Ҩ"��^Q%��Hw?�g�ݎ�1F��^�A�����C���J�=`�f�i�x�)]h�CX�;�C��<�E���6�|�N��j��Kc�����s�W�l'��%��Ր���r.okFq����/&D.��P�$q����ꅞ\*YW�4O���Lv��h�Cj�m�3�(��p�R�H�%r6�� f�ut	/Wt�5��GZ�m+����O'���O}Aok��V�!��N#��gdî�������2�ÛQ&�1!O��4�.*�r�y�ܾGQ��6 $������w��,?8)F@1�ыZԛq��+���7��U��/�~o�8�s���WӸiJ�!�e� ���8�߀S���̪���kp�� `�1C��V�7����w�7�=�3�;}P^1������t�
��;�J]Rn�!)u�9"�0��L ��@P�nA_��.�	�� �6�
=d}�St�
Ϳ������ ���y7K��Z5��.��W���;Ȳ<��xz���בw=���� 9Y¼)�Xc�8��5Ze�f#�aS�OψuQk��j�w���4�ԉ�@#X��}#�v�Ns����%S\!�?t�"��A^��X5��7���cp��01��p�NZ-&�j�+ �B\�k��N���K���B�xs5M�[cDA��؍2�4(&"�ci.'�=���w�}+�v}PM��]�Z|q�M�1'#�ܿ��NC3t�#�w�$���dX�RA��ȥ~��h�һ��g�%?Ra'd)DH!s[���C�Q�<�GU�K�	JB����Y%��,,1�O@��q���x�A�7C z�fl�r���1&�_�r�an���g�T�fq��,�:��g�4D����vq)�>�RC)f8}v� ���rg~�j_=���
��*�����$�{̔'Rc�U륕Р�r�`�D�71_�� �K&l@Y���`f�����{_�Y��A�>��&!iF�R	����)�"BʕպP�B�Lb��}�lM���״1�<�E�s��GE��5�7O�"b�!�C���M��Y�5�6Z0�:�;�Q���O�maş�Xi)� �r��q���C���S�S�!�%������TjYF�O��3�?��u0�G�����T�(�ӑ&����ȣ�K����Q���-���-�XgE �{F0n�X=��Q3A�Ak�� Ad�{
�$�ݶza6�)��/�S��;�(>��M�������0�S�����@Y��m����rZhY�%?�@<Olb�`���~�m�S˜�4v�ԉm5D�l�0lϐ<�*g�#T?�Pk��i�n��4��U��2$!		��V{8� ��Y�N{P�ex,�u��BvK�w�����L����3��u�M�f��E5��ߊT3�dy��F�fo�"�(��wd�e���A�([� h��)��X4n������+M!�7rEH��Z�>wZ�CC�ƙW�@��R�;Z����M<�d�8��ci\U7�S=�	��Lq�4��霄:�	Qd�U>/�e���Qh篰/�ٴܞ_G���{�T
\���V�уV��v�ZtT�W� lm{�"�M'��ܝj�H��>�j�,"k�sY�;Zv�c˘��nj9#���	��:-}BN.ʓ'-4`��沂@-"�3��`&j���kŵ���$r��&	˨�U����h����&s�������D���A���N���}L�)4�T%T�R���D��6�1ؙ�4a.�����/-��b�:�Z�%��2�
:�St6���C`{��I>�:�̎wjwL��2T ��r���k�x����i]�*���T�~�	��:�ws���������⽋��y��)z��8m?�M==@�zU���a�����f(8^+D��-
�K����E�"��7Q��> .|���˯����n҃�7.Ts���X4o��H!������Ѷ;��R!�j���o�Ȝ�_���P�����c>.+{�r�,k��θy�	��?�� S�_A���dU�G�;'_"	�&l�.L/�L��[!MVt�üc�����h�pżt^�?�.�`XB,ǅuD0XA�����+Z��4�&s�)�ׇ��j�H��s�1�㥧K�)w�b���-��#)h0I��?[P�^��� �F$��ռ�?,X.>#G6�HS�#2]�U�莍8��wv�j���V.��|�=�9�tq�{�
"��9uV�5#��M��׳O_&4	#U��b�4C���Sus���O�\N_�
�ٰ���t�'���~��l�m�g�����b���b�|
��ֱ�?hv0�_����C�=9�y��Yʹ����篪��1(:/��qߎD�*�;а�ѝ�G�����+��o�t��)W�F((����xn��?.��S��;W�B�2�+� 34��$��pA��m�FJ4H�����u��yi�l��fX�e�`C
�k�S����Pk�����#@�~C����	�Kj#�w�3a�eV�v3�|Ju��+�0��J��J�K�f8����WaDmGHQ
�������/�B��uڷ]n���'�Ϧ���G4��f�7�w` �Q���@��%Ҏ+�B.�V��Mn�'_�BO?;������h����R4L6��߼{���I^_�_�M-Y�:���N|�r;X<�D	ns�w��4�o��@3� ~���M���v����/�3� M�Fj�w/L�Y�pgBu����+�$��TU|�(DǠ���/�F�g-[klV�rmc�[ե�k����S���<H��=~t�'��
����e�:߬�8P�cs�g폪�#Mf�^T��y��y3�"O0����1C�����b�,���2E�Q� �0_Z#�N��O�L��-��,M��=�<A����J�Q�H�b� ��Q��P@��˰����ԣ]([�N�T�w��eX��}�Z���0�^�OP�%6*���8\��3����Y��,Դ3�w[+F����ك�_��=Θ��C?߃���n����%S���2E���j�ޣs�X!���6u�p��a��e�M��w��mG��<yî9�t����� �@a	`I/\��s�I�9`d/]��^:���ݘ����O����������+"��/TS��0&%w&��thv�\.�ySfUykaԖ�0�ȧ�J�����h��¸XQ��TAi���9��Gy�5>�����u�S���
�h|��ES��9�4���3..�!��+熂�LLx�{_u�����~�1Z�|�WI��~r���M�.��G�l/ �p܉�mk�R�gˇ�}�%spOF��4��rM4�i�f�΅��2�)뻖�W��9��E����x����J'�2+�h;grp�α�vF4��uWW�:.�Z&�ѐ������L�W,K�CC�NZ/Ѯ,,����8,�~�/��c��F�=�|���7�A��� �{f��f5o�փ��P ,Mu�Sk��58Q�Ⱦ�)7n�:����i��N�����[� ������Ae��������r+H��C�a[)a1oT78g��(U:P�� S
�MUq@rq����a���W�߭���*y��y~�9��n�M�"�iW���#՛�Ŝ�h���L%�H�v�}!�ܑ�	
��`7�7���I�O @�9�������\�iH�{	t�k�]MV2L0��}�Ǒ�	T������{��JN��3�&���7�y��Dv���q�?7')�]sE3��o�ɿƭ�9�ҿ��CФ�OLz襁O^X���q�[�p��m?}@#�:xyS`&�w�)�oʀw�[%�)�{��<@fqW�bқ�d�U<���Skcv�,���X{���Uk�����Uef���$��L�_Qw�顂w�vܭ01>��e��u����Y�YR=5��< �X��iݗ��m�WO�����q��'� C-�����r�7�_�*e�����T�*B�0#=��%Wp����k�Q.;�g�}���3�%��Af�x�n!?�ɱ�!��X)3}����]��n"��v��I�s�O���lד��EV�ӝ>1�U-9�9�F���8l^�S��ʚ�9�l�<��~�Z��_�Z%���U!�=�����`%�+��B�ګ�#F��l��6M.K�IЅ \y@i�(���}-+�_��͑駿�J]�\E�<!n���.g���Ԡ�~��~�ض7-�$���ݼ ����	<�1��O+�F��oa�ơ�����f�!��>N�w��^�P	>�$�g�����"s3�ZN�0��d[�Kx7+��m�O����������*Ȕ�Oo��.}��{�������P������v/�)�ʥ=2oj�v���PW�^) �)��]]��9���]��;��*�!��� ����iw�Y'�#b�OK}Z�YV�c���LU��A�!dR?|
YvF�ʫ���1ZIl�"p�7����y�!M�љ�2���ԗ��f��P���������ݍ_\ȧA>����B�Dlf(��; Bןj>�"d�7���J�-����ͫн�ʐ^H��pQ����<T`���*n���8���)]�J�r�i:^�s^��h�6��0� eh�AZ>{�-�췁"�#���`��O[���"c��	�Y��%r�.E�Hݼ&�0�uR��Tt,�8���^
R"\�h[�l�5>>s��~����w�u�05��m֓'��%�����v{��Xj�Yܥ%`�%CK��?���E|��]��98![b��u��ULs-�`2Bi4�x5w`�����Â��o����F����t��\�}�5����7���0���������t#����{��*���tt�]�,��Ȗ����11����
t>��w�U�����}̆ޖ��Ί�I�+��>�7t˩V��8_�{ʶ�B}���c�nѩ Д9���⺀�ϺX�r�kvQI�K���_׻����:{T����P|�z{AX���r%�$�23�y���}n� ��hw�����_Z�ǈ�^�#l�;�lQ+���+G�U��Y�r���C�ΐ������i9�SƆw\~��d�-�r���<��� ����7Ra1T�Ρ������=��9����L�鄤2�Ϭ�4i�Hd�b�P������{��*FI����m��b��( ����@����8��;a{bl��`5�$��xZ���r��+.�h26j������~h�ʩB��ҥ����I�1�ɒ�j�����-���qKL�nf�ߍq�TԚޏ=�<$g��ٴԴ^�-Վ�N(�h�5����(^x�����`β�@~9�L�?�/2��d�	�:�QFy!@���OoLy�]�B�D�u�K~[��FDy��#��}�D��~|X9����L�)���NٲoN�&��>�/P{Ad�"+�ʋ3��@]��}�����ū� ����b���gXt���i,���u�:_R�c>���g=�_� �G�M�֘f��V��PJ��}�����d�<��L<��>T������,�اe�Ҿ� :�#g!K��~�לigym;[6M��ʜ]/���l[ie�9霨^����x�,t M�=��P �p��Dg������)�'$����c����d�5��'�V�-[{��4����c���1rMEO�W#σ�ti�T�1�c�c�G���\zI=�1׵X�QN:�s=��w��@������tz5��\^�ꋊ0RQ�]��KY|����3T�j���g��;��w�m��1?W�����+A���p���%�3�Ï3��Iٍ�4`�ꠍ78_h�����b4fl�JZ��cX���T����vD%d��jkc\��=hs��5������F�PF��=��oR�ǬC�k	:e�#��PlÐ�@/���8D4J�ǚ�N�/���^P��l=1�pKq!��5�2`�G�U���ڦ0�ڧ�Ϝ�2�p�dBG5��'L�ةj/v�vT�5�#��5շ����g�����"_́�QDf������M�hA]����Yg�filc�v�,�PD*&o�ȁ{��d� GZ�˲DFk��lpN�6%`�Xtb�B���1ש@�aR�kpR�:F'�w��%jR@��G��!���çr�1Un�0z �2��g0/?�X*�A�����u�E��p��&��,��H)u!�$![��,��Y�M��o�7���)t�-��a�!� � �^�-���l�ɞ�8I���x�1���±��Ro���W������X��\C�<���i�>0���7��*��^�[�Nb��w��^�Y�)�h[(�u�P�@_A{y������V�WT�����A~��E����H"2��uA<^��׬D�0�yӷ�17��h�c�m���K�6�M�p��g��)lڇv�^ �^��l�4����7a���m�? ����Z��i��+& ���w�ùP�Z<�7ZP��W=Q9LiLY즫���_�֔i��/]OU�hv��aSh_T�"�.ap�Mms�>1�
^#V#A�վv��p���B���S�fT�%2-V�����;��h4r�=y�0qw�X��@ ��s�ˡʕ�X8���ޭT���]�9�����Q�����M䨢ahf���"ו��L�u�� ���1B��O��?�L��Ks_乹�TH���#tk��S��6Y��倥!�R�:�l�E�N�`�#�x%����Q�����E��ٿx+�?���i�p�=�fA_}�h������0�U{�Ĭ��ݩY��יM>h��^�ْ|�h� %�3�l��Կ���*P��J~�<a�"�Ozy����wk��p���`Yq}��O�$�Q���J��(��e6�.с����zi��v�^�����D�^)B���lCѲ�����m�a�lv��{	^��Ӷ����Sq߷l���P�Z��%�#���54	@�b�5��Wh�W�+���>]vhܼFM���rү�|ښ��0�68��F>zN��E3t���G�X�!Ն�k �z^KԖ��<�L,GK��vN�9���
��jӖ
��jq��/��g���g��k�~�sqD<� ��ͪKE��%Ί���5�V��0��uoVB|�`/��+6�@�g���΁�\�k���vs�]���"����e(��eR��Ou��� �4�<M/Ri���Tf&2���s�V?]:�bn��`���W����rP�8ܧ^��y���R�&���,UpH�cV��7�'l��)���i\N�VlqF+�Q�Rgb�0�R��R(�N�GX��}Q�o�NT��a�?R<Z��B693��E�i}�΂����^OR���|�N5c�|D�?%0B������)������0���6l�:���O����,/��V
o6J̏9c8�F�Q>���&!s�����\J� _��XYHDݡ�3��[C�Du1n|�����Y�;D���Ē^-Ԟܔ�T<��M�LE�[J4����b�!'fh�4�xZ����%R�n�¸��ck�Ԧ��bm��n�Gυ/eD�[�e�R���|/>�A��Y��};Nr7K��-�k��k�遠D̡��op� ��t&��
������72����Lr��0�$S`��V��<���?;��L�b��>*!�����D�!F���ˊ������
��	�Mf7����eRE�,�
~a�`Wo���.�Џ�9��D�g��	�x,<�IVZU�c��b��J酱��r��cSZQtd���}i-;u)HF%�v8�hX�B�t1����V�Tm*���8��ĕʲ5c�%6�4Xbɸɒሏ�0��A+J��Qc���'��p��p�}��S��ߨ���F(,J ���IQ��?� �$����)4��k���
h��Ju���^,cO�bW
�с�іv�A�۫�Nںwz(p�$��w4�!/P�)-��qEvYUm���=��tl5��k9x�PrB� Zb?"��*f���$��.L��%D" 7�<��D�m��X�z�,]���&���+2bp�R�L|����Ue��/��!�Ӑ�����E�
ӎo6�g=I�H��)-�Z�֞�MQ�3�ci�Qd}�|�1 m�v$y���~K��,���z�ѫ���\g�*��*E�����'�
�H�w׼ag,�;���,�?��L1oxly<T	�݃��9~����bD�v[�T��A�a�(qn�� ��a�ʶ�N�`��"��XL�u����j������- 8�>���V�O��J��H�`���������M�R
�Z�9�H��(�e��ۓ�ߋq�?^�=$x�����v6��U&���y+~1z�G��=1��<+�k5C���"�ka��#I�)fef�z���������ۍ����l!�X�s���{������5�óH��p��G Ɗh�D���)*�@$܃Id�!��6�;�;9jsYAu�ޣBd��5Z	�WD�{7��釕D����ت�r�.�E��k��5���y���{i�G����ĝt��]�5��EP��r[�P���(��ķ��˃푾��%#��VcW�"�@�hsl~�c;)_��ɇ�>���˞�G��[[��ʏ����qM*�� +0;�e��/0�G2�\?c�!>���N�(��=��[hW�;�p��Â�B�5��{�+|����H�Rv���r�&���'�O�y	y�|y��ǃU߹�>���l���*s>.N�	��8�A�|w� �tt�b���!!�"��/3�]��ĆԮu���I�5$'${H}��8A1��؂}� \~y�ţΊ��o��m6��A��@��s��
/�R�8��as{5��w7w9sȪ��1�HN��Ԑ�o�$��a�KL�O����W�<3��1�/s ��ᜤ����J�j�E�˲ )�����K�����W*p����׵D��]���!ϻ>-�V��1��Xa�~�^*�R �P�3vXrrm��]��校�p������YŜ�l��h^��j
+�l��j���+��ێ�d中�_+3O�2v��A;��.Oy*�g��9vL
����Q���畯���ZP�����(�D��o��wn��ڐ(I��ߙcs�~�/J�����B<»�7���
, 
P���B�\�p��K���=Un24�C$S�F9�R�B��iE�|B�Ol4JԡS��P��L��P���[�0TO���u��XZnV�d����,w��v�B"�K,'I����PmKŧ�*VU�����.�;�p\�E�s��;B��n
�Pc)����	�7��=h����CM���&�~ȶ(� ��}�� �[��e�q����1˄��'��,�*F�1�=���Bғfc]0M�UBn���V�א��=g�$��*<]Rg^ 
�ɲ�ε@���kĀ	´��B��@�'�?�����y���~��`½����$e�tˊ�iuiEf{n��ҝ{��?��d�J�S_"�k�_�)����:�Æu�)C���n$�t:B�,��]����md�I9~KO�B8���V].��`7���
T���gEJ��W�)C��Ԉ>��n�ux$%�$�Ю�M:�dE$:�L-�b�<&ƌҕbw3o��D:��w~����=Zy�[�(Bk���+˽�X� 	F��bf���'��b=��aC�����ĕ=�Sd�ӭ���g�P_��-�q��@�Ƣ���}u�>:]f�k�`�y5�4��*��z�Cx�����< �И��[�];�������l����K��a��~���춛�K@��=$���$�xl���wEy���_������|���b��x-=�'n�R̭"9�*�2�~��]��#��^��������p��3���e:��(���__��%����t�� 6��ه&�=.}��oI����4WiUc�ά�\����=��?k��3O�E^��N9 ���h�T�>��:S���VL;�c�y�!�]K��e�p�m���x1T�Q=�i�!��I;s�-���K��5i1xgG���#���@ˏ]z�h�.<� �������y�j��rA�+g?�^\a�;�ğ,���y�6��s3�k=���e�Zs���R-x� ���^I�#��c(P.+��>�X����lG�V^(_�C�ΡnK��>C:V���)�(��,��M�5C]JJ��J`N�K��M(5j	Ͽ�ev_L>��ӴAÃBX47q�/�y֍<љ�����O�|�M|�Z�ڡlgH����j��s:�����0U�Q���t>�R)zM1�m4U���znA������tg��*?ݚ�2�D%ƈ�U�sKw"r�����'ʿ���Y���� Zǹ�{u���>�Ru���-[&�Q�K�~�ڗ�"׆qb%M�����������m�-v*n$d�����|�"&�A����5��7Ł���{s�g��A�Lć�/U~��wq�G�9�}�}ǝZFʝj���f��u�Ӝ�����n̩�����Q�0���=<�d9W@aP��|�\d｠���wSA�2�#^JM��hDo�s��$��Y�ǋ�	�k�/��j������q.E�]]�qc���w�����1�S|Q]�yJf1&>X��5�:0U�
p�?vv�$��	A��n�0z��5}�0�:�aM�'�� �2n
�w�г�\b�n}�Se�󌔖�GJ�7�4itCZ�/�e��JXM�������HA0A�55��<̩��(��*�T/�9���l�GY3�����G��tJ��A��������y���g�ā)L��·$g�%f�>(eټ�uxH�����τ�v�K�8b���*�/�����!����~�m��������o S�Bi�h����Q�#4,c�ɏn��O�a��1+��gO�=����][�yV;�"+��I��z��Oz{�m";V�;x� ��F �{��8$���p��gk�4�6{��Bp*>ٰ�}�
�3�GgZg�s��������qJ]�}�X�-[ Pz��� V(����t⯙�tk��Ꞙ#���e4��o��J!IH6,-�E.���0���k�z}��d���vWK���?��^lS��^~�D
'Q��gEi�x�ڔg�VK8��ژU��e
6_����Z�7�J�g���hkU%��������ɾ�/��r�N��6�t��09��B�D�������|kN�7 �/��2��bh��	�!IO=�4��[47q��ňA%Pk�aOw�3!ǂ��q��:��'��EX�ɮ6�ق��dxEzJZkTJ��8L�z [�qrWQ2�vU�@��](�,�
8���	wQZE� �׊����b޸��
ʴ��������[����-M��Q�uf�ƭ�@��:������������u1��PM�����zCZ���1@fx���:$��X��R�č��T6���u���א)}���akC��4%�A��v�t����7��CO�$��HEv~ۿ�پ3c%_\# t� d�r�BY�����{jl��>��� �{���'/_�^�<`S� �"��MX�;�+�Ų�=�>�M��0�!�|���8���{�O�/�:N���ɐ�k��g���U�k@ _��1�]GԈx����� �v��}�zM�(�=�y���]�kR��
�2�����P�7���&(-��ëY��̴춵��L���v�K(�t�V�R\��q4V�=�g�z
��F!�2s鶂��I�(;��7�4ڦm���%��16������7��rg�K��F }Fډ?��D/̽��k�b��+�7+�\�J.;&9T^v}���^o��窟E�v$�(]:ۍB�.� ����'j̎�X0oW��f,�[ս���#GF�������Lvu�W��6ٲ/2�R4'�
B+s+)���cZ@�����E�ܪPn�N�ڞ�ٌ���2=��N���� ���gAX�~��MVt���e��]�n��`'P���#x��ٸX�J�Gr���O�.�)���d�����"H쯳��%������`Nq��U���ەké��U)IԀ��sԿ��ݕ�(��j<�;�h2���^��� ��a��?��i�[nLWC�d�5,Q�k���T���f�]\��7�/�!)����[��<���(\R���)/�Oxp� /^{�,�u�.ա�44r��g��H�����e�IE����K(��I�
�zZ� h�Y�]`_�X�2|���seyp�"N������{�jˣ`�tg�1���mF ˊ���-���ѩS@��qr+���&�i���T~��6B�gX�s�s�ܱe�`�[�#�/���Q� lܪM9e�:6��7��[��B� ��&�������@.u>ɉܩ�����"N%�}I�c4�MM�#qr�/�b.��,�[�'��b�6������
-U�V&����@�>�h���B�N[��'�>|�Qxd.y|�8�?F�O��w.�ɨ��?�P���}O�t�r���+֤�G����g`ޥ�rUj����bl�ϥe�E��1��Lq�PڈB0�o�t��ԙ�kU�B�(��3_�g����{�"����5�<���L�g- ����4�s_M|��B���L�	�Kݦ'��w~{S�4Z�! -��ݓ)�v���ƏքW+47�g��fB|�#��g��� Ĳ�� T> (���M٭TcY)�ٿ��vW�f����U4.�#z�&��hv�,%�+�+�+�`Rc���40��p&�������fw��� T��;�pF�2�u}�G`vo3b��1���e_Jh�R�������y�?�%�ܲ���.��=kC�~
~%~*�t�k��ӄ~*�RRR�<6� �)�������������+�R�K������T�h�l�R��/?E����h1�՝:� �U�����LڋPUm�����}��>�����]�I�b�čXC��Z�x�M0�Z
#��V��?2g'peU�������W���s�5��|�7)Vz����j�9��MR(�H2`�T9?�Z�E�4�.���
��T�����Kz>y�,���ym=$il;�߹-����"�%.Ɇ��p�Yi��~/��_K��|����7mtES�V���*	o�Ưΰ'�Z��b(FJ���&7��x�n�l���+����q�D��Ywo���k_UN]������`VSꎀ�7%k��b627�(�ɠ ���-�^����7E�/������\9j�eV��[�.���p��7�֕��j52�H�u� �H���fҚ8!����Ύm4�[VGZ�$��@nj�Z�m0�MP�$z6!0�����r<���e���g��J��#��O�� ]<%���^Vߢa{�$ȅ�����d�ɿ�<=4��.xF
��VJ�%z����,Iޚ������y/l�'w���`L�b(dI�'��?j.�q
̙�LL����s٘����V�|��$��H.��P�!e2 v�T璘a�Txi�uC�>��3���R7��fD5@�j<F�ѡ�x��rL�|�2ޓ��UW���~������7]�(۠�78��Oq,�i�[������ӱ���1	􆓥�̽^�X�:���*��;�r��г�W��^(��!��Ys
�hD��u:��"�9��M����Ϡv��Q�;���/�[��+��&�5�T��u�F�+f1��fo�+ a]S7O��T+�D��w�D��"m��'89���|��?9,�d�( �/O.�8Kc�â*&_R�����X�|��7�ޏ4a��gF��u�?O]Vv��9�aη� 8�dD����2�M ~������L�\ͫ�4Y)g�48��8b&�F~�U�ڞ��Z�#|����!��Ǜ@����\e���!X81���@D �i����B�u����7��8!QQi���UC� �<װ��C��eB���^�gI�$a
i׍��ݲ&��&<��(Wa�H����s�� 㕿C��ip��e5�&�] �4�9��?9Y��E�.��N�y��A��J	�t>�f���3�m�,Ft$3Z&��n���+��f�kb�B��rM4��"��鍸e�v�i��`�m�LV��Q��k���E�l"���,A�U)�D&r�Gp2�ڦHi��7l��|h16��ukտGb)l:Y��_PB��(tANV�^>L�;�B��`w�6���?����,���r������b��]r�T%z�0�M%�{��SA�V6Ғ��1+B�D�ڜ������%֝5�/v%�����,lt�b��T�g�`������6GM	��}��/.N(?�{�x/N��d���I9�|Lh}�TM��]���ZY��E�-�0nkW�٧+[Y������j-�E�?��}��m�,.��`����؟]P1q�G5&-��F��^9��Z��NS�ڣ)��q�C����>�s�h��ƪ��O7�_*���%J?��[��p��E	W1R=�'���R���ِ]��E�����G���xxӔ���9Jk�#�O�����G�v0Yly��ܽ7��.����î(I?�&��ܜ�����}�t\�T�DLC�QI�;*��n�mfyS2�<���d���8�Z6�6�l�A�/3b�_{IF��'_�y'���[<��v��kEϋ��&�����(�����i
U��*��r(���tU�A=����� 	�^oz�k���mn�&���o��e�jq�����
�X�Uj�ѱy�H�~AxaN�dz�p˅3녁�MBys�Δr��3�q/fLk5���&K���QL�L�j�B}�3M�\޷^N��f>���[��'@[�[�\���� .�>��8�G�,"^qA�f�R��ty�ъ��y�y��xWiҥ1_�<��4:⿓n&譡��-�?�`m=炢8G��7��U����������1��7� ���>Rk�y,����Sc����(�Ⱥ��W�}~�-����p�R�f� J�թ�g�IIj�K������������XyyX��_63E-�:�A��=r�xB�a:����o;�{����n�
��)<"^d���YN�r,�@Kt~�7��+$�`�7%H��̢/"	B���&��4~_�A��N���*�vH�IdD7c�?��^���V+��͍:.�<�+����̕�ZYklGȐ)�{}m�P_%��9�J�6|`e��an�VA��1=��9�c}5�ZZ�P�0�U�2Q x�X�9�v�bW���p�a��
.��a[~�S��ٯq�dpq������;c%0r�I�"E�J�0^���z9.V���:*Q�	X����h�R�ؓ~�44xc�����t ��5C~R�P{��?r,���2��}���(9*C��� �}/FȆ���|�e+�*�,�H�z�y(�2�H+�
g4J�.�-tn�Y8����i(Q~�K^��#�(�B�t���6���$��X́�Gy'6�<:�-��3�Ƴ؍��j/�0��m���hR9�����B^��%��S���v�N�Byn'J0�[�B�f N��hiSj܋-�4�G�[�ǭ�kW�WwƼM�8� &|�����a�2ݽ�{[f��(ގ/CF�?+`J�DY=""�.Q��}�!/?�\�D�����k9�
bD^	�#���:�Ah�,��^O)������?m �Q�?��ĄN�4�ԮLP,��VP{�%{�P�pZ����m��1p��qM��&Ga근���oDi9��-!�����f��Xu��qO�7�3
ޓy�Sy�b*���B.A�o�������cP|7��g���B.�W��"t�#5��P�N��������a^�͊l_�_d�Q5�ۄ�� #����q���������7���j��V���<W�V��I����M�~��Z��y�Bif<�W2��⥑��@�et`"J����9]��`��K��#�Xe蚜�!+��1�It�=�6M�k�C#�bǟh�R<~�b!3oDG�g.ꆹ����3��S�}:Y@s����ML���#�hʍǁ�Hϗ'<1L�}��=m8P�.��}$�yn�Y�b
vV��H�G`��B\��D���f�#�kt�� �����E1!9_�,V[���Ǯ�ۛ�a��65���;j���±^Q�ȫ@��!��(�����ƝU�%�q��ۧb�PO��y�"ygI���.�+6J�0��ZL�/�+�\jg�	�6��?�9d�6��v2�z�
�7�u�[�c�$����H���<<�}�"b��X�.�ۑ�$�S6Ÿ�e'��ԔW�Z�ֲz�GNt��8>���J�ڀM�����y֬bw	�=|��+	�UB���J�k��0^�����D��.�LN�1�/[YF��!��Gx�G܍1i��~[�+E�ֹ�ᥦm�z\�)j��(�y� i�C<���ϋ����@]��Q�FmB;�4���m �$���w���%���Lۑ��_�������~*Ԛ��)�X�kO�ϞW'�H�l��)�]6��;@u�]��;fR#���<n<�{��Č1��Я�5K-}	:ϛ�����*~N�C�0�lĪ���(��T����;xät�BUW����ҶT���j!�8��A�Y=��I?�=�R@�����[,�S���P�sQ�ͬ�sM����qFD��(5��x������*$��>ͳ˃9<R�����!���hS�f�\|2�e^��Ij�N47�W/�+I���/܌��t�������Z2P�̴��$C�k���|e�g�)��y>>�
�����f���������	-h��k�e�[��������T�0�\r��ۢ�>�3����C"Fw��R�6LC5�6P	�L2����CQM��"�DP����T���-��n�`(�Ȗ2|y�n�L��'g'JV�x�D�Bv�7��B�p�hQeqM�bO�Ge��4%R��L����ׄ�!�����ހ��y���V�&��_���t$����<�����n7�Dc#�A4(��f�-���ܰ �_eG.�J�0��/`��&��(f����o��;��LA��*�}�?~�����e4$t��k	EWJ��
�Ike
(��l��+�촴ݎ��GOH2g�t?k�b�F�v�6�p~���_嗅���!�z���1 ���`�k�xZ'x�bX���H�����4{���4���8��z�O�z���\e�g�� m�@� ^]�G`�&���Z��b���zUB>DHl>���н~��θeL|>�p�)۽!R؃�6�:?đ�7Զ�c�u���8ga�uY�sx'U�Xex���1&5���HO��in ��g�%��sW��tn��a���I��
i�E.�H���Şg~�a���폺kǅ�S���PP�*��_�HrU�-�ͬA��a|�T��YWJ�� ������EG��(�o�Tz��Կ��>���oVbe�����h$�`��6�O��:��6�6ԑ��?��5ٍ8�ṣ�pSd�B'#�c�D�K�s�����7�U�9�{*�:RF�D�Z7�*��DB1c�^��/_��y�����>����Hv5\k�J�U�aS���L�"�݊l5�?{tQ��w!N�lg9}ҕ�C��am�%#ސ�����Pf�����R�k��{l�D�3 �ZE&Kߐa�ս�a�V(K�'����x��v�ǃ�r���g�W�&y��4|V�OuDq��^������L��I�������9�'�	�Ϡ#е���3'_y$��*��(�����	r�+���E<Bj�\;���ڃ�U:�}��%��~e>uȣk���|fF�g�Dr��U��/od����e��R��B�f��|�,���H4ٗ�z��ي��p�J��A[�U����Ƙuy�P�o,׈�T��4�����9��d���-m,�'�\-��2�
�����vu�Ҋ~~���-���k����b���j��ᚌ|jr=k��7v6Ȼt���~ɚ�fC��
7����	�)�����ۗUU�q�j����+8N!�S/Mu�F��:A4����B_.�\��hR;$�0���x��	4��8�cӘ���w�nA�V	bPn���)�h2��qv�iL�&�t���P�Po1�~���)_�}5�pBj�Җ�_ˬ�O������31�OϷ���w;�T{�����>4)��J�Q	B��{������ht�j9�)���W��Fq��~/0w�k���z�(L���p�c֖D��~C���]��Z�DU"6��V�D�,J�>uWj��Z[w�Ǹ3'���kխ	Ը����MQ��/f����bH��k����Ñu3Q*4Q*�&P�M���Lm,>���'�ڰؼk1�ā�p�;P�����V�'��j�b�����n͊x>!�N֌��άO��ľ�:x�ʆ4�)�􊼋���Iӏz@�X�~��Դð�cfv;/���f�$;��ŭPR1���tL�i+����h>�pg4�Scܙ˓��(woKi��<�R��NQ�_R�����P����.�j�{�M&�����c��$��@NM�1v�J�K. �q��[\{�g4F�����b�A��7D�c+�m)`?� ��
�Ǻ���@�$e��1�R�Ku��[	�����<������˅!�*dOǾ"b5�M��$�c�f�Q��<����1�1�խ�o&̏�a� _�K��"ݮ��Oﵷ��XRϻ�<�Ɓċ�r�io��Lr�[2����ț��ʫc���uG�K���k�AW�e��=�<`_&�F�eү�M�P�cg�
�$����x�iBC���Ql6�׃�(rQ�@`�x����_|���0A.m鹿`g��gP�d��d5ԡؐ�"��/��L��%,HL����N�C�rr���t�/���s�E��x�"���W&֐���J��lX��l�?K�=2�?������x�'���ص��AFV>��P,��9q��xЭd�E��k��o�8&)��wڎ@��X󨅭H���]���u�J��9ĔV �l5���yZ�y܀��P�{A0���s=�e�OvIy���%��#��WY��� �w�3l�rO�y��R�<�S�i�(��M[f��v�Π�ilbmm=(R�ו�c�G��l��F��n/M�D
��W��I3���gA#�,��Vt"*��L��� )T'5,���՟���m�Ǝm�j,�û�Q�5@`j*'rU��%��s_�\]�0R:�s��3�~s�<����U����-6 �GWق\��듯ySŎ�^KQ�Ę��P�t��عZD㻏:Υ�4�r���U�ʉ���F�,�j�!�C��w�iB����� �rG��q�����,�m�{YuobN�`U|��
�v1]�^NgJ8����l��Ѝ$��_$m�I��n$s�x����F���Qj��-}c>ʬ�vǞ�cS1��"�`�������(�℮*n�@�T����5`>�q��=~Y�|3�O5�Sd���d�����.���-���DW��\�)����	l��͘R�2��x00�}m��v!�;�A:/ж+}��sQMr�琫8W&�&��p�8ݦ�=3�^Va��y�X����E/Ԯ����T�;�<��Ͷ���h�h�4 MG �UX��:�'EM�Uʠ(���� �;"7�*��&Z+�Δ렇�����W������?�w��DPpUC}e/p�Q��&���дo�X%��3!�b�Q��ɋQ�!�JFX x�1m���� E�\3&ؘ�J<Ř�� �ס�� ���0� �f)�r������KT�\��6�O*�W�omǄe^_7��/��yJ�0~�|H���ޑ5�1�p�,���G���>�b�N[Z1�IC�!|lI���=;��c���%�"��Y�cU�w�R^u��������T?��P5X�֥Fz�Y�x� L�Q;N��∺��}��v�];p�̉�A+g4DL�K4C��4�-pʌ|:R{_t�����h̨�z��/2�PIhϭl��u��:e_��LA@i��\�򠅷�ΔèZ9�"ȃ+�C�6�|2Yk�k�A6ᒂ#�9���1��=�s�ᅸ��Į���*S�A[w,� on뮞���[_z}���/�w�]ˀ{�)Dz�m�Xu���ǫ3�����a/"f)�ǗkřYøM�x��S��ՙ|���K�������Q|Z�BΎu�>lm�
�pH��l�W� �����D��lW�H�@3��
���P,t���@�N�`�a6�T�Alg�4u��L�݊���6���v�0%�u䗘�e+�F�U��� 0�����I��Wn�M����p���io�fL���/��r�/C�:��r��+�O�� �B�hɝ�B�+���.� �߈f�=A��w
;�k�i	xed�rD�%�[�k[Y�q���&��;_d4��S���p�籐wu��j�fu8wb����H(I�t�s�W�lͩ��%x�� ޷�;�+ؗ��w���T����e�3��xo��/?�"��Ek�����NW�� ��`�mS������Ա�H��Ծ֮�R�E�_*o�9�u���|�z�o�,������tl�j���u��JlQ�0XFu�����'����=�]���saF��9�M����wy�7ކ7�f���l�B.� ǚ��Gn~���pA��խZM��SP��y_f$�) Me�B�s�6?@����I����)��k�T,��9��(O�?�؉�qb�3'�+���J�3�<D.�)<q�l���E����̤�{	'&��_}��+Z!9ʲb�iz:��筑(rL��z��d�=d�ɏ�Y�b�n�]�V�����pc��+AmG#D��(*.�_�qg��Y���ѿ��癅QX�(��S��O� l��Wz����f�dH�s|��8P�8�M��F����P9�E2���aC��M�\}?�bpհ�xj_7��pQ��{��9��\Ch��F���Y%"~���)H�~�-�Gs������c�Î�${S�?f�k�������9�ơ���� (�D�x)���ڣ�K4�
ɝ�������f�9�?r��_B7�{V��,�����ن��k��k�pd�����U/�+V��G������af�wD�F�å�al��Y�D��2D0�ď՟-'�;a�k��^�ŀ����!��s����6���#�Ǔ���HFk�|�I�����7����H*C/�
[s�:�.�5Z��ID"�[0�X^׽Դx���{��1T��룙�:�t�]���r
r�����A���M�r�bT�^�b���!)'.?�C�P�u�+#���
��eG",)!�p�.�T�^�SN�m�a�:��e �9�6^��&�3 Q^�+�~�V�w���N�V�$��:w��I���S�`���f��!�:v�W�+���$59������$ܬ�� �M�m[��Y-=1�T�u�k�@�lF����SR�쌘��}S,ϳ�N\���{C��DYozv�᧶�Ξ�M�;nw*�k)�.�ˋ��x!h΅�DvJ��a���Nql[���H�$�]e7D�;҈м�rΥ���G���*�[`�2+���� &� �����A�F���{I��˱��>RZ����y��x���*Qm�^
Z�'�tm�jIO�a�귴y�'���T��#
�OU(��
����*{��;�@�j���2���$�`����YY�I���w��s��u-�v�:�54���ŵT���-X��|��ŋh�`����2�;I�����f���Ae�~n����hQ���6��������hx��G�&{~�)�ɜ�U��`Q��y�<@e<Ƕ���6�q�#�2�K�_�w�^��� ���.��:� E��tF���qYY6i���Y'vG��=�<H^�z8�n��ϝ�.p�jq���:OE���B݇s�Lhh�Aߔg䭑G�8q�%sip���\���g��.D�c�<v��j9���2���79�d��.�`�:x��|N�&
������!�a�~�cL����΍;/���<X��(�0I���<�h����n�c�1���o�q�2wBH".Go"��h_�����-X@�\��.m�p� �TG�8� �aU{��n-�!������p���4�fGgd.	~&zi����� �m�۱��?]�T~�y�I	?)z����(���#uP6cb5x�{L̷��Q(ݱ�h�P��S0�`��H�+�8�Y��H�Gc\�h�-8۷�h�v�S�2�M�Jǃ`���E�G������j���h>�8��|,�j�|�lM�WM+F�b�}^ne��}�'��'��ǧ����!�|�S��T�~?��O���K8���%b-r_�����g�?eC�(�*_F���s�/[�׶k*ӮW	G���BX������q�UVz7��O���)3�%���P&	j�7[[��z
l2�HdN�ڄݷ��`-�8G�)3Ղ�+�s(C��w��&�À�TYԛEA��[�wml9�1�a�Y3�G��&^?�ƒ"f�Q��`ܴ{N�D֬.��4���ә_g��iXB�G����2 ���{�7p4x6�$�"���H�z�@f�>�\
��ǰ۵�?\.��W����*6�K��B�8ºu��@�'�o�uG���~���}��i=S>Y�`1R�#$�Q�҂�J���[�E��F;�i�\.`k�X/���f�k����tP:�=�	(LW
P�mp��qt،��[� "�B����cYPl��A�-����<dh^�7�{GC�y(Ѳ��_��>hZ��|�P)!,�q���(?��~�
�W�o�/����#��6L�C���<6������+>�
����@D��1BHH�T�d[��������b9�h�Qw��M5���t+��:�'�k�E��z[�\��V�⶙1r�H�����1���-O�	�ll�Ɯ���3��'�ψ����%<�P��2� ��&)"��$-
�V޽Onp-��)GR\)/�7n��b뿃>Ԯ�Z8�u9/Jh^������J@C�����W'rf�v�Y�w��&mgn� �����]*�4ld�}M��(�Լ,��!d�r&�+��>���*4W��0'7��˽�1
�ۖ��8<!T��A����q�H�����r�3�r�˾��/����/��~���O�Ϊ\�\c��`�M}b�n$$������+ ! xq
�6Mߔh����<4@�S�o�Jϔ8[�o�p����t���K��a�n�ˣN�G͎���|�"b�g�e������k�ʙّ ��\��n% ���T����sr�=�����ܣ;|��S�����&1"����?Nb�.���s��}��������XdT�]NV��Z�E���8 ��}��z�{�����9d��g�[���:�k���c���_��OH5	��>-�n�]\Eii�x�B��aAƳ�Y�D��b�L��f���Fݫ:��u!�u�DdH5cd,�}��Z�*�Ё���+��,�<zܾC�+-���ݺ&5.�h�@m�¶优�Bw��|p+��޽��"w˲�a�n�a��� ^����{�+T�#q�.�Κ{�)�^�~\ ����j���c�Q�
,q'4Ӷy]�Ur��Y���&_"T�߫�CC��mh~��׼�D�G���u�,��9�􄒴���]�*����nG�o�J?�M�eyELi�k�6�[��ӟd���Y���n�eܕ�p��9�G��n���)����4��ژZO1�8t�FW�b͂"��h��>:�Un��zGkK���K�It�k �EQ�bHc���U�ב�d����]`�e���L�O~��ּ�r���V�}�:��,��jl|�6H"Gt�VP�cuo�oz����mT	��F�j�(�v��M���^-�^:���_%t>�nm��~�0�)����/���PVJ�W���Ay�c[(/�A��.�xN@*W��}g̽;�t�p(�
���;��l���R�`%��Y�5���O��`|���S|y7�5x%�p m��3�_���� 4sa������4��
o@��}�%���ǐ�s�r�@���b�7	�4�h�>����q���3�*	��P����FR�o%kf��| A�r<4.��^D�!�Y&E2�G�ՙ+w�ݍ�dN�_�0���j*GE@�7�ڮ�(s#c۳��w��Q��NRx��E�d�-򇛓�y�Di��d@W�ſ� �ԑ}���Iqm��)'	U͗�Q|�F���]	P�j޽�o��
a���2,��=J���2o'�k�a��O�[t�r��N?����ʇ�08���_�۷�f� a���x������p�9ꥐ1k��	G�	8�3�W�J`U�r�Y� Y���w�	H���ߓ{���!
�F^/��^�8�9���u(? ԎN�!���ݼgu?�0�B�X~�Z�Pg®��MD�#J������Ul�:�@�t��v!�9��36?�֕���l.4���ElS��ĻJ�U+5N���Y9�E�s^O��A���*[�����X����v���;���#��0fW���i�u���6w֒4a�z�r�C�� ���Xe�a��3r��m]Y���*&ϱA��D�W����hx\?`�ѭj:f�G֩m讵��A�+˭�������j�<8+}:v�i�S�@�=�����cN��i�;���u�y.�%�_�8G(vb�7�
��1^>)��~�:|Kk;wG�@b���p=�k2X滻IǎJ���\pw�M.��=�=���dU~��xP|��:���V bE{���w�����>�Y�;w砉]��h�P�B7������9�i�9ֽ��W��vZR�����U-�-kg��l��kh:���ȝ�-�:��� \�n^���6|R��Q�N6N���QФ4��}��{\A��4']���z`��Q� w2O��}��
�:b��fs�JF	HE���Ó#qP/1����u�J�������P�2���.b7��"��y����
zϼoc0�Y��|��6���7�V�_�}0U�vc�
�S�LJ
G;�*��am@D+/��n�������B�A���x�a.s��s��	��1����������9�\Bs�T�>�3����v�C��i��G�8~��:���J\�2ld\21�[O�[���7��P���wE�4��f�P��e&���v�_Y�x�MvN��%y��s�3Q������t ��6�P���t����k9+]��V���mC��6y���Y
j@AxZ0D���^u"w\�x'`R/4��a �ĸ'b�lg�D0�_�ċ�%`�/��p��k_��9��C4���(�Ǣ�%Xu���f�8���x�S�u��!�	G��@��Yu�����_��Q큺�ܜ�_+/AGn�bO$Qw~;�E�]'�t���IH�)5�[b��r�,�f�:�ED �晎�Vz���k֗S!���΋��<�h&��h$��� }k��}��Sئ�.�_��E�`:;lѕd�P�u����	n�Z����[�6���2��i�M\0O�O���N�waN�'$�x�>ņ_$H�rX"W�'��^r�x��?�,���m��:O�&&�:���.?�۰��]�v��&Q�ǥǚ���_2�^.���5>�sT&l�<v�����Uv��{�0
�a��'@�mJ��ΙQBs
��S���Q��� &�XOO)8JQ�X��A��1��C}U@4�M�k{�O<3Z�N[���O����zaSѺ`�J3Z�)��g���靪4��$V�6g���Y���1V�I�=`��6�̘ + ���v���jWX�;'M
��T{��x�l�8^���X��oP��l��&pD�ϰ)�9��L<�J)���-��,���|3�� ���!Vqj�3���)V������ԋ�uIc� \�N�V��Te��O_� lT����Y�����~�@A`	B\��O�����e4K_ڠf�8���X�	b������N��R:����~���T��#��|���Ə*৳K��ɘ�u�~��Y7��IՔ�Ýa-y�D)��@��:�0��{N�g�d�"0.b�&���@́(�C��`�|,
��T�����l ��	��M�^�G�����]���S���F��ڋ0����u�%z���<	mۚ��zu����BA���a�?6�Jϣ��2�^��^���z������	��QӠG a�m��z��,my���.�D���g9��"J7��2�b2-U��q���|>U�?�y�K�݀�o�>$	��V#��H�Y���w�d����(.�CA��a�ΘI-�w��BJ��������#d@�Ҋ`�%��*��dv�|c�X�)"'<|x�[جo��%F�
!��xw!X2�p˼vģ�Q^m�qխ-p\�$N�I�A'd~T��S�Nr�Â�n�)<9�?�HD��v/>`�.?#�p��J*=b�����P�u��ɭ��,s/4"NEQ�
�5��_�<0�P��'R��3��.�C�s򼺜�W1V����tx�U3yǘ#li��E� �H�~s�1Z�@����I��%T\΍�l�������E[T4��I��s��RDq�֚��
~�����-���[�3Lq{�ѻ"N�lj��	��{㈯�B�̒��Aw]8q�ǵ����ɸ(I0��s�1=|���]u���M���X���/����m��!%��dq��:��#̔Fs�Hh.���	�x��!�����ߤ9�)���Vv���р�uÎ�b���l.7��h���A���I
I�
���)'�#-ƚx��B��ׄ��?K>��1U̲Y�b\�n��H��R$F	���g�\��U%8u~��;�'��7;=-H��K¿IA֧�K��T��B(�Zs*�z���c��4��晱$g�~�T��z�d�N��e��xΥ�G�g>��g���(� p�x��/Y �RD��ڃ�;"�F�>W���tƆ��k��ψ�Yy$��������>�n�m����b��{!��G�e*ۂ�7�O�U	>�i�eeL��-��s��I��z��z�/��C'��T_��m�[������b0� �>�u����S��..��^��k�����=�Z^�����)��{��?��f����B)u�HJD�~E�A�;���r[n�_H��u��-��r?�þ��T�5/4߶^��c<i�����T6),#N�5�C6�4rR��'4��L��	8��e�ȏ�3JΉ��e����B�u�"�d�jk!/-,EbF�=�js:q2��#0��l�#��z�����j�5��Qq;��Wѧ�*}�����VO&���>J[��2"���)]��u�P�9��SsA�|$
~����5��i��?~g���l-�Lhf���~�&�������fC������uݢ�NT��W~�޺����3�
�YD�
�=�� D���K��ކo�3�����ى�f�AdVS���K�)c�i�(�a�I����}����6����׌�pL��A�����	�3\p��A�#D��a?w���]������s��Bw~D!��^�Up�h+��q�lc�T����FA�K�";�R~Α�[:�e�eM��N��ϕ6J�Y	�)`�=��B�0�R��{+m�p�.����8׊(��$Z��E)��L %�l�ln�|8�E���^�c<�5�����a� g9�A�>�C+��u���z����W�O"�u�B������K�&ܑ��mܝ�x����𘦧���h��`��:�"�UCv0L��u ���y�^E������¥Q,�C�*�C8x��B��۵�ÇUM���j��Rtݿ�u���O=y-��q�gy]�'�xu�-c�I�}��c��&?�a�ߕJ��k�g������NW*#'���&�mp$�*ꊏ�܊�C�?��Z'2�����O�	��	IZٗFxx��®��h�Z���E��Dޞ��xG���J)���[��?Ɖ������O�"���l�������{S���A�㫽Ξ&�Br�<.1gX+�nZ�8/�:v��5�X%/��s�����}F��� �0
���������B���N��XE?C�0}|}$!����рfKu�3~=�J�'L� �]�P�v�ur��s���JA�� ��%B���S�P�W �x�+Դ�._�eG����A}�0�hy��6�N��ġQ�'�6�+>v��p�{c�˷��\��,*E��^[������zXs�`��ʤ#�$�$�H��*^j��WV��&ů!>��LH]�_:�s)�gν�\� 7�rx:�<��_�!�Sڌ(97���/ >c�=y���z��F"���6�D=r�9yuv,�1��^kD�bv�l�1]-u�y�_���t7'}ޤ�uJ��Z<��w��y�ޟ�R���P@5��3aZ�sB��=& ��DL \ty-]`f���L-�I�rU�1SW�e��&,����7�W�k㈭|�K��O���Ÿ�С�:�2�<lh���5�h��:�ه�N����-��g���{o���p�^�͈��)g�`�Ot/)�w����mo�k6�;�.Ң�(WO{4_j�m�y��B����O�4Lmo��bn� Z}���9�=���!_y��M�L*
��[�VJ��|:�u]�9)���t��Z��)�/��J���qN�:̵�q��R�%�܃r՝��QߘO�nu�
A���f���>�1���f^�&����_ \����9��f�,��ē(0%�N	���<n��G���M-�B΍�K,.�V��N����s��CS�hO�Տ��'�l3hU+�$��w��B|�nb|��δ-Qg�I���k��N���_d٣�*���o��3��@������-���(��G�_�(���,_�T�"5���ri��].��f���\�!0��O<i݁�,���{<L58��'r5U�sr���b ��?U�`�� Jm��|��7�X�����n�D�ʳj-^�e4���� �&��T�{�=0c��
�I��Io?�O����4��,W(��~���6a~צ���f�Ǳq]�HcJ{f��	���O� pM� \D+k��F�z�ڴ�QN��Kc��;��^[������פ�VU�:_�zO��U�pL�GVi����������"�\��@2��hD�9%�������%�7h���녦@�2��DT���{1Og��!�[Y#�Rݯ޷���G�:=�-ڌȫw0�bs�0-Rm���U�d�y
��:DB`�����*�H�t�Ǔ�i��fXj�"�.��Ɛ;^s��-tdC�3~��o�*����-�8��b�g�$&]7 �c�����b��^�g��i�xl�(��M�5KQ^Ê��e�݌A���ѯ�]7��S�광m��"ľ�b���U�f�ې��]�.�<ƹ7��~������1��*\PX��XA|+"kHa�1u:�Q��f'>R���ߎ������n,h,`xϙ(j��G��^�rM����)2k�j��<�����@�al�zj�9+C�\\^Xؕ��/��c1�1��ڄ6$2%��x �]�}��-����}�ȿt�JZ͝�9yX�Y�����,�g��.�Ҕ:Pw����^����E�}$������J��rR�停v�/��5�0D�����{�	�*OC�k��,BX��" �����6I�D�B
�H�0b�m�<����������b;�&)�:1���]!�U�E��I�RB���#!�X�vf����P�����;ig@8ʡ�*.\|p��3��#����U A����B<y�m����J�;fF��BbEtM��naQy�ɚ���R� *�M��;3�,iv�|��X�G_�r����v1��	u+d'�AiCz_��a
ob��1�����;��%�6�
r \�aY��_
a�+k�1�����B��@�鑂B�$D���W/��m�? �k#�~z(���]�9�T�n̷wM�a�� ܖ_��W��2�ܿb�_��x���!5�#ߚ�pbd�:�|a��*˷ �G~C���T�`{!��7DYa�h�����q<o�mLn�EM�\=�-)���ݽ�\y��Ybc�: k-�8=�K9��ٲ�u�}z��l���	c�G)h���B��x�ץ/{lf�\�#NЁ`����1���<��W�����ri��D�E��n�A4�2�u>#	����ԙJ9�&����vgD��*���2�6�(?�f�:aL��y^�X����_SRګf��@	Y?�!�.���ɏ�����}1�P��Ul�!݋"��c<+94|{���z1�<3�<j0A�Qc s)�E�{n-�s���^�T+���GkW��@�NB��^�E[��=t��4=��c
B��VX�#{��uN����6�����B^���_e띐�
�xiv�)�䳼�������QL���8����^����|���������Jm0(4�犠D؋�d�;����I˟��7L˗����dP�O��&���k@
�d�k�n�]�<�M~���ۨ��ۖF�I���-��9~(�|.�����t9�x�^��cM�ُ�o��.bT�1�>�#�)��F�N���������b���2*�L.�Eh��,��.��oTΔ'.m����e���|��KH�g�3{. ��dY�0k��⵹g�����9=-�FPe��2����O6v#���=��՛3w[I>��{8��c��	�lP��������ał�u�ͼ0TƊ�/�<�����-o5������6����02x��C񳘋&y1�"�W=�$�i��������~�b�� �x�ɷN;Skx�Z�o����H]:��x��� OEK0��4j�q/$w-�� [G���D�2�}S��8S�L�`o2����Ō`���u��J��2�_��=�ay0 wE]�у`�r��Råݷp@��E~5M�Ŋw��A����ʃP���D��>�Y�lj{�dSҜ/�?R)X �=�?���'a�[.����4nV`�_s�\>��&����sP� Eb��8�$��wf	`�O]�W�dR_���ޙ)>��tՀ�������ϡD�9��x��ܖ��>?*,F�U)5�S���}�R��c$X/*����q��c�>����S�5�Zl�xW�U�= zU����K�Ӭ@�T�G�c2��Z�Y$�'\�Ӣ��C�
�K~g���ݐT*p��zG�2/2~���b�&N֭��P�:�8�	�e�E|z(Y8��o���`i�pͭoČrQ(���\Pku��ȳ�B�O&c��݄�L�5��>c��>�1��
���S��̏#g���Ey�q�{�;�b�&w:�G����Y���	�7�QDP5���1��O��L�1�J}n�Y�������aO=1�j'V�o45����!<>�k;��4>��F��ܶ�k0��s���A�S��"n��b�~��c.��$'5����w-8ω4�臞ž�>���w�j�~���Lb����r'6[���|j��ذg7���{���ۛ�a{2�y����'��>���\�߄'U^#�Yk8�ɵu]�a=�8?�FQW4�AW�H�����ll|� �A [��]���=���m�x��,�!���`|X%Ŗ��}��i�v�)��c���7���e}ҳa���t��
Մi�Li^ ��˂d$u����݁i����xJ����MlC���Σ��d�ʹ�<
3�>eP�Xm��O�t~�?�}*j鬩��2��tIJ��d$���pG!��l�e�d���o=�ie�-�gƤ./��#2J�+���,"Go���Xp�<h��)�D3�]�_���/@$�9�;�	����I���}��h���
}��
�N,a�\_Ry���X�;xy�8��)
�m���~%�2Op�V��U@���q�7�'ym������k���^���h[����(G�3�����O���LZD������V�>$,j�� �Yb��������<��SKfg?3!f�����#ǎ���T�}��(�f�'�ꪙ�{?�"ɮ>�t��`�+��(���=��Hqw�OlB��nZT�g��Ă.�fIE�Д��o����E}_м�ީ9���9�2'�Xm��f�d�H8��sUE0t�F��_ˆ
�4/�v� ���<F��^����;;�B�;��h� D��P�GK*�)�S�����%�-7`X������,�!"@�.I#5��ja`uf��J��N�أϑ��0�i�,������R�a�ʼu��;�yb����������ʙ� sd�?���TŖO<��n_��4���1[��_����]�\�lK�z���9�(ϩ}.Xt���V����F�9����H�?��&����f4�
��:JX�Kï �K��n�rK��*��M�$Es����	�+q`��1cB���E�u]o�*Q�%�`
��0�|< ��8�����{��FO�0s4��N��:Ix�g�}�>�^9y�_V�:]�>5�������I֤V���2.񌱈�]��~!4�f�Di�PQq\�=>�G�Yz����'V(%acg
���hغ��K"UjO�N���S�F�%�T>��Zn?���n+��N�<Y�R-n7��ۼ�N����P�g���b	�x�ڼ<n�C�Y3����uI;��o$dQm�2y�� b-5�K��J���4 �q��1 A�-�T.+ͅ�X�e0 �lA��ך����ˊ֢�v�����Ɔ�ќU��?	Ne2�kugb���l��ص,��$�x������g�E�%�� ���Y�<�.���;��/��n����-�!��ֿ3Q�淁!�_�4J�u��c�B��k�U-�tC�Ⱥ'H�G~aCq�U��g=�6T�;UK_���8mF'6����p�j6|�R��1��Ꝑa ��gW�-���_:�(9}F�(�?�"�q �.�����y�fF�h�HhK�	�����a���25�O.�_VT������dyN��^��{�<|�Af�|0lt`G^?{���	0�J�N�o!/�/��j���	���h�3�$2�p�Z��Z��ט� ��i�0{��u�~�7��]��l��(��'#�m^�	x|l�n+(�L3ؔ	�e@X�¿� ��X�O��Ta�џ��ƛ�;�R%<���K�p��s��-Q�`J~QE]M���8Bb�N��a�������`�|���M�9�����^2���������q�vn����>�R{}T���U0����
�IB�:�������1ᜟ86\[���Pf_�
C�+9?iJxA��5����d���K�_�E��\�8���X݋��VN���\g�◫h�R�jx�6��u�v~�J���i� � ��/�ç��{ůW;}N#$��Yۜ�y���=�mĺ|��=y�����a�
�T��R@4�P�5�(;L�TW'f�;�^HyR��z\�w)x`�a91#��|.�-(�MF�;��y��6�Yi~�k18c5��fo�ߙFI���G���./1��P�D~",nh�g���"���f?����t��Ȕq�$�rD�|Y+���U_����1����T�T%�]���c)��0��.HaT�����D�`��DN��hں��Ŀ�}fr���1�%j�]�Oa��1����M�I�'�U�k%�es���r��.��(�&�&����ħ:���
	�!�;Bk�|GOQT��n�O�T��2�N투v3¦��;ּ-nE�굈�b�E��>_l�g�Li
¼�`e����z��<�1���J,�/��q�H�x����*����v��e� �q� A
:�d�"b-���U�M%Ɓ�������*��TE���k�9����Y廘`(!Y������NW��j��>���Zo��g�g�.�,V=��l��N���0hS)���]m��-�:�ֱ_5%��웏؆+W�:@��������Gr)aʒ'ɢ<�5�s�w�IV%�y��B�D��?A`"��u�(��l�x��!'o&�2G��|�=r�ǟ�ȣ_; "�ww8�a���u����BH��;d�SdjW�v���?���s.V�@�hӿ�A2O�`�"T��(w�1��6A&��`� Y��q�t�&gF%�̷n���g|�rw��P49o5UO��F�����m���%byc���� �5�b���ޅ�a� ���;�L)��T�M�K�����	%l�o�g�{��l���m	'�Rn�~K��0��(�ʱ�o@H������n�Mٟ��ho�\�7#'�y����#�8�)�"�������9�:K�nIP�1�x+!�\��g<�A��V#5
�V^[,U��K�	����0�T��+C.�P�'9N����9����ʖ�&$���f���e'�V�싂*�B�P3q���b��[�Ly��Ā��d�$���ڸ�-�������X]K\r��%�2�q��[��|�# ;d9(e˶A5�g�F8�q	��[�Ea����a�u3�I÷c��|�d ��>vr_yl�)H	z��J�mj/�=)����G�L�$�La�G�B���+Eo�V����	n�Ͻp��ʨ 5��D����N@5���qS0�F����g~Ϲ���.9j9��	�`�� ��7S�I0:�S�hc�䟱[,��Ӫ�0q���Pq!�0PL48�Vlm��J�@%��SkSw��G�Zq�|�t�!�9sYjj�cX�qEY*��V�ۜ	�#@F"��k�p�Tƥ�A�G�
_�򊆅 �5E�����*���x���<�Ԉ�N�= �soT̹��q|�&�_~��N�?�(�:{'�2���z7� և�8�B�4p�w��a{[������l��F�l0%���u�O<v-��� +d����8C	*�5O�����ZوK��0UN�_l.K�-�>b!�!VL�=������No�B�t��\d�����P�XӘ<��B�!��N�2���9������F=�|�'���d�e�	生�3A��J���;`\�����N/\��/�M��fI�̞��Ҽl�Q4b�8t������y��dV��7��,��9���Y��ͦ��\W��#ß�bGJZ!�an�f=,̵���:��lYΉ:�H��QX1���Yk�]��Hw��Ǽ��IO+�L�����Ҏ��m&SD����t�����.l����&�?W|��Y�h��e9�)�
Z�S
�p�Q�.o����פ��13|�2�oҙvYj�<B� R�T�|�*^�j�h��݌�P�R�/�G:��y�d�x�f����tIU��<�s:K#w�����l���/�i�aChL9Y�Ƕ�L�=�$��m�^��r�(�i|M8��F��d��FO0Y.�Ry�[��1OF�׫#��Y�{�Hkc�m❪-}/�ˌ����)���L��S!�"_��ܢs��.���_��Uv��P��u9ok8�Ň�/������>l=����6�Q�CA���r�uiFm�bS�Q�>��$������z��i��k
�Ƒ��Τ����Ԛ	X��G��c�U� ��m�����oom�+gpHH +u�>�9�G�"|N^��8�)`M<;ou�Ӄa���;��;��w���WJ��k��ڏ�\p�<飽HG��?����e���uu�l40��~�
�H�v�Ef@1С��|U�{[��1��?s�Nw���K���(nf�X�j��]U�G9\	m���?o�H�S��7��Q�{Bh�@���Ro)�pŦS�D�Д>&�^��yʽ)٢����k�z�ŮD���4��B��b���Ҍw}e\�aF�^�X�/��?�ҕ
į���O#X�I�d渑��/�}.�S�Yj���,�wH'7���1@�Y�,��Fl8�]�FZ�fFs���o�V��W|v0���R8WE�^���Yl�ad�l)�^��1���z�yo����� ���j�Ƒ<]x�Xt�s�_�8���c�Z>�Y�5A��Ӊ��	�+�� �����;�����K�l&�GA�,tD����"�I�@�i���0�4ID~S���zBOl��U��+��Ksb�LQ����^�S%��ϋ/���ϓ�<P�٘�Nm&Rd�-���>��u���-"�Q<�����;�.	�n#������Z^.{�K�<�/��������0{� F������8��@��m�U4�E�/m}���A7d�GN��)k����8�w�#|@р��U�^��Rߴ�2"%�[�o���+ejϰwFy8T���dtSa�xh�s��h%;��*l8�a<�%dx�'�{쉵��Y����r�^��G�GE0(Ʀ��CU�+(z>��6щKkԱ�k��y����?��
,r[��U ��>8_����h�!��U�
�G�!�59=c��B!D�A�|�md�B�	�V��������|�U��H/?� �����4.Y/�j�
�[�v?�n>�z �7$K��v���[���S��[�Y�����Nۇ��\��I�^A>��M��1M�2+)"��e4�� �߼I���(�X
l��!%iܣ(��O���π鏐'c.�~���A�]*~���8Rx4���� ���܎vC�� Wȫ[b�����r�
�}(�}eU�@.�	>�A��A���ϭ�p�U�q��{V?Da�%'~x|�ԩ��@g�@��4D�١c�@����\3�W�퓳�����6�*������>�������%�;L��J�!�����ZF�{P��I�i�Z���+=*��+I�{��U$�?�%���־Ua��X1T��YX&�+tug'��ɵ¹ȅ�_#b4�%�~s�FƮA��	(@�sчPa9ʌ�1�$$�����n�-G�f�Ѽ��Z��Q��),{�`�\�ӈ�ߥȔ��&ޯ�Ȼx\�)Ĕ�d[����N���&�z�sq$�t������QY�!y�HQ�H�_j��?κ��(�5UԢ�2�|g�ta_�:H���aS���*�uk<A���������P���C��>/�䕛C�رj���1��d� �v�3"7�T��k �mt	�rC��v[F-�k�����B��T{�����営j@�2��M5��9�L&���Ң��V��J�)�*97�ࡓ�BjҪ�P���eu��r8 rH�E�ؠ��?�������Hd<P���!Fjy��};�p����mG��3Rl6\}#+E���ΏF�LN�!D�3w�'oOM�{���m�������z�x�
<��]����k�V7���0����	�ب�&N�l|+�o�>����g�񛥎�/ "�+ic&'�/��x}�AZ ao}>R�>�a�e��F�]��f:�d�a0r���O���z68_S}����y�1�x���j�Z,͇V\��|`��Ւr��ۡ�NK29+Re�*�4U�җ�¤؋���)��+֡� a���t��I?Wm��O���A��]�G��;�$Az�7�~C�\���2
i!��NV_��"r�f ��$�ӆ�чu�	�ܠ~���=�s�[FHm�6�V�E���}��(��[���'w�bdD��JM���$�Ñ����'ڝ��K�)Ji�K�� px'Gh��`��R���b"���z(��I��C�^R�7=^d����G`�2���vSk��cioC*���\⤴��-V��W�qe ����F�8�hn�UG2O�BE���K�&	w�# ��:��3#D���0��K��U����Ŷa����6ږ���qҺWV��o|�ߓ[�y1�M�-t�2���=3U��]��x5=�iim�9]��h�[���1��k�g��@�+?M8��stg<�L"��	�'z���w3�;Mm8bU�)ůEaI 3lo�2�k>'����-U�m�f��3�m��=A>Sa&��Ǆ�8G')�Wf�%|qa��s��|NC��L\]6�hL=� 2v|b��M3:c������w��n�e���6�t8Ꭸ��;�XA���bG���ߦ	X���ni0�(�����\� F�W�Ko&�&=Xp�ρ2���$�pXoE��;͐�LX�8��D^��Z�&}��j�u2c�(���׫-��[��tסW�F�ܱ�#�ԋq�$sP<���ɦ[�K[�}�H��(�y�T�|!.�K�����*��#H����:uJ��*$a�M�L�|dR��*$Ɏ-��S4�U?���J*t&P���"�[zC� G��z�^Ej3�ѩ�`���n�ύ�m4�N�0Q/��)uDs����ld&�U���خ�}����Y���$Ʃ���q_<e�P��NC5��־!�C1�Tc� =n]�p�֤WY����:q�"�@��5Ӿ�^���p�t�c�by������5f���e�� -	;����pY����X�=�R`���`OwO�.E�_����p��ڏ� ��D�vJg핮�^GXm#�^uC���}�qp��BD�z�Kc���l&�UG��/q
��2�L���IQ74/��H�8\5�F�"﮺o!��Ȉ!�.}|8��ݨ�r�`�2���%��?��ʆ}׏�O�qh�ct� ��=����A&	��>x<J�QU�`
U9���/�O� 	߅B�"�Ȱ���0�l��3%�TK��l�Bk��@��r����{)�-��rQ�q���ּ���r�T~�d-zp3�����z�PA��bw�)��n?��mg<s1R���g�ho��F��� ��Hk R�������[�<�x�<XQk��H��vB�m�oo_�]_wL�q_��M�9IxK�@P d��]p�׻�ݦ��/�q�d� �-����Ҋ ���>f��`J@;����Zeׇ&[_����W�����̽G��+%OC�5e���Ý�5A�����m�����$� 0�R�'x���y���p�{�a1"1����Rr�l����H������ƻ���I\�1�i�Cc�,��5�ӂ�W�\b��U˴��yx��Q����=��#$�������[�$��>��w:p��Z�k��^}�l$�wę�S2����m%Oϰ&�P��i2ٝ>!矃��w��V���]X���sC"���J{�6 X)�+v�ؚ
��V˾k��vRE"y�?ۜY����s3��&Ee|�J�rM�@��(�LM�H��s��t�?"g��>�)Hu4HNνC���|�]<>)�'�Wa~@�w�>V�1	��Ba�xF���	�įȖ�*�����+�&����*������
x���P��[�Ex��c$�e~�>���-�F����U��~�������C/1��f<�����C�:dɇ�]Z�a�O�(Z��kU����������9 [@㙅���ᘔr.�$zq�.�ORCH&hH�4�Ի\�D1�*�~��VX���Eʘ��E@���B:!�6��|z�~��%\Ve��7O���j��g%���P��w��U�S�!�������Ϻc��h��L��M��da��Y��͗ �n���ήux�N�*�g��;RT���qXm���� W?�� 0ָ�u�%�����
1��e*ʢUx� Y�a�ɮ��hk�Adcl�kkĜ���J��
���5��4s"��%��
�� �A
�f�c1��!<��o>�[�O�)�ov@�F��Z���U/�.KJ;j���9��=���?4Ғ캆TE�����M��tZ��Z�Wruٮ$4k�?25Qm�Ird�JAA��?�a07L��G�0�ֱj$xj�N��t:r�c�J&��|�͖~�a9Q�;A�B2�a�E���,~vΩSD��~��0g��$-�
���%e��A�
x���<Q��B{
(dB!ȝ����C:@��紨��j|y�G�5����T��؏?%��̶� �����k&��G<0jn�ޡ^}��MJo¯	�H0ѹ{`TnrS��}� 8����ĐS�-�t��M��x�_0�?=���Z+�6�I륲�l��K����̷Pb9�V�lǌ��Od}D�aܩ�x?���̣Xc�M��%͏����qO�G��|���ŝ��C;\�gFIy��]G�*\��ѩJ6����������nR���}�n��F���2
q�`�'�c�3�(z&�����J��\^�� wV$a&��aW7B�:+�<E�ES��.F,A�~O�(J����ӱA"�V�a��q���!���N�;E��ҏ�̄�A��4�}6���h�vG|���/r��@��"�F������T۳���Q6Ϩ_T�O�\�-��;�	�1Z�,<��h����I���ۇL�h1K}�87 ���]�����>�U�a��a�mSz�n�bg�� ������x�
�����<E6���v�KES9P��} Th��S��[�o�U����`�e��)h�'�x���'�Ӹd#�vO&'���V
.xvB��eZ�L��Ϯ����:�_��}�C٘���?+3��R������!�O��g���i�V�a��[����.�@A%8�CT���.=F��� P�XW��<���c��mH
���S�����◾e7�����ҥF�5"2gJ��4�nT,+c�n��e@��p4�FD^�T�BS4���;���Z�2�0a�^�\���k֐��EP�a`' ��`�]��- 4�Q��H'�S,���ZK�6 ��q�=1����Px�s6$º-ظ��ke�@�OxQ�T������Wk��w�J�1�&��03c�Q��v���Fk~�ǭ�@x���4(;3Gb�kݹښhތk�W�����)[]յ	�x������p7�J�
�8�24,�d+(M��Ǹ�<�	 2�8E�U"��n-^}Ҝo�����:��>�7fpEU*7�o��J����v;��sOW0���'u_P��7c6����l�Za���;����[�d�X^�?���
�"�� g��ċ�Q���QH��I��IH�^�;d|����<P��9X��0}3d�Mj���@��I�uu�51_y��&<�o���*|�l��ժ|e��5F����]���,|���)^wn�v�����5Z�k��߻
 ���>k�bGC�v�2�v[D{k�47(�m��lkVĎRX#���pz7"�bﲍ��	���RσCJ�:)O}�,��P��?�Y��bviI4�EFy���������y'�Z���	ZI���Hew���3�'��3ݖ)�@C��==�#gQ��s��7c�9���Y|����������>AH��}���Y�"�噕W����S�������gD���L�!���R�L>�
B�yy����)�N��q�Yp��?F�b߲xD�H5��
0I]��O����C�Χ�T���(O���O+�:�[�ڙ=�T-�T1�h�.�g���"�-X0�,�� p�Υe@wl'��g`"��4�t��X �Xݱ�T$5>g$�Oפ�#����e�-R�t��@~��xت����X��O�i?.���c�v�����`P6�`��ƭ"٦�r�����G���2�6'`yM��N"�,�<����8Z�ݟZ	A#k9`�&��x��jj��+4FAXB7�f��!��Fif�wIT8;�W�>�&�H�@���`~��$���3ώ��_�Lݠ���KgQ�Nȱ�:�2�g�>{��N`�H�q޽�Bj1[��-2׾���A�M�}Պs� ���=]��T�
��[޾B��r�g�6^^#�v����`_y��:�^�+��1��(l�2�=]
6�b��?v��Z�F���Z<C�$�����S �O8E+�3&CN��e[�k ��V��Þ������ނ,��:��ׇ�bΚ����d�� 8�Ͱ�6��*�8� ����%�|�����4M�*34��R��%d*�hN ����P���oɪ>-l�z�bi���&\{l����_�J_~���z_�5e�$m�z1��`O�f4~��agYyh� 2oRc��c|5��Ǐr4��dZ
��=��Ț�H��epJ��i��'.�P�~??mM�⅖�()�U�s�����>�M#f�qR����I��3���y�s�2v��ټl������0V"���-�Z�W!B�d\_��!�k��S�ʸ)n�|V�񅣱�*��f����"^�P������a��X�B��U�@���įz{�!���ɴb�Y���Ä��`	����_�U�qW��R�?��z퇭��;�Z�� .}��[9v}��!X.��-�C�@�_���M8������r\���p�8(��sQJz�c`T\~3�!2��ѪDp#�zY� ����۬]p�f�/@�;�+Ź7��u����?B�Tj�f��uga�M�Y7&�)�C���IȞ��EOKC�:fi7,T�4�4�E�-�.������0?1�/�C{���~e����)e��G?���Ɵؿᑥ�y�u�Au嬫z�ٓc��(�~��:0̏`U�Cfp(Q�H��g��텗�J4t6l��4���x��D]��?;���n��0))a���)p1T�G�Q5 �ф{&P�r�T���"X�e���s�k*;ЎO��,ʅoŠv�k������u��4�˴���������;J�\q���c:�A���څ�X�1�^Ĭ�g��&�j��[vO�3���{�svhB |�rT½�C%)�����w"�jн�at��BO�f��?l�K���z��
��<�±W�3��O��l�}�4��I�4d��2kW������ڱ�ɑv²g,�W[���o�Z]P2k��|ٮ���}���crw�ͯ���IԔF'�ET�ƨ`������4kۈzI`W;�i	�!�U�)�8�˔�;�����šO��#O���L�2t#�q}e����W�\	.L�:E�����'���v�`�o���� ���R��4��A�<&�M�z��2]��OuF�Y/�.��i^{��tH0��d��h27�P�M���!V�*���0
�-��;R_�5!�i'�
 �0[���*a8%6���c���������NVn@i���<��A*HT\�)�����	�2e�'�z<ߚ�Z��E��6�EYҭ7P����>z���tC��d��L8�0��J5 P��s�F{�ʞ ��:����a�>��I��9���Dkmj�eќL�Ull�MI��zDjX�s��S���4���y�5�!-��ѨSߛ�`����6Y�R�;�i�;����m��E`�v�;P��yV�z[�Ic�sGӬf�A�������(Ș�֏��e�����9O�a>���)f�%,=S�G@9xpU�S�4Q$�)M��+y�m8�W��
m�R�|��z
UK��V�qd�_o�1�����'���괋���٢`,g�Ξ3H+H۩9`�+�z�XnV!ժѹϫ�'[O�֎�*䦘T�i�[!�[�2��jM���p	�#IgGqOku�,ߒ�䆮�\�yV���X�տp6����!�Q�Jۅ��F���y}KsD�B�h�7�䠨Q��c+9@�ڢ���R1�e6���7�AJ�>?�}�v�"��L#��1��|󖥳8�b#ZL;�{�B�S^:�W�Ú{�W��N�cA����w��m|�bn�[�x�:��b_P-R���%>L�_�����+�_Ƙe���%R^�:%7՜zt�� h[Z�	�p��L2H�y���~kFh��|{(}�F��U'ܞ4��_�>Z�!:�͒ԑ�N'���V��IW�<gs|F��GD(��c>{�3T�F����a�>c�b4��X�o0+3*7��3�#`Hs���D���J��/£�=y�a�C[�����w�n $�w�Ξ�=MǴr�P������g�:�oB����8�.�d��\wx�.dj�f��U���  F���Ҷ����4F��q�������)\���3���.�� ���Aʂ)�qB0�uy�h�]/ww[��;j��%Q�zxD)UY���^R8�Y�+) g�.�l|X����G�'�ʌ?I�yC��Gώ�R�6^� �Z-���{F�Нs��&$�_�(���)!c��g�{� K"�x0����{�=��W��V�tڸV��.�rM�@:�؛�ҽE�W�e!_ZX=�Q���0�7�g�=W�o`.���u�.�i�\��b�F�V���Ȯm��`�x�
}�
��V���|�������<���N�#��L��7�]֕����%�Y 5���09
9\:�8x�*�������x��^��3��D�����4r���$��&e��b"��P�q�)����@Aj����Ag��&@!��;��q4Ƴ�?�ٕ;i�d�?����]����W>T��Y�M��َ���^�[���0���T���W�!�׷}U5�����zĜ>>�:�����H���mǁ�Va�p���D9���l�s��	�}����GD���?Kz��k]����|��"͹yCv	+̈U�.�|�0�}��J
�`���/r;���]"O�d 1�i6J�^c����)�y�������Q?C�(���G�Ҵ/7�v r\�T�@�c��	U�����W!��)h.)�ӏQ�%_��Y��|���SR�0��̾Nl�J��������#[B#��4$�IF���U���B*�������e�RN)�it\~J�Ƕ,w��=�#�H�/#�����T��Cᒺ|i%�S!�Yڕr�� ���P�{���Y�p�����C�tM�Y�����R�u�
���ʷ�@@#]S���wTt��>%���!#v�&�O�Aܦ'&�DQ�;&w�g��W�������d ��5!����zm�&�(a�"��I��_m�/�z��m�y�_A��$���ֺ+͉�k���'I�R�f,U|�O�G
�	����!�ީ��d��;�!����S���i>67�����S'���- ���(��|'d�~i��Qg�4�T�-���2�Щ�=���p�/*���.�dl����V�	��@���{��Ltp�1�Idy,m
v�)g�,N���Y)"{���j#S$�Gҽ�X]!��<�w���D�҅x*N�����VHރ���@
{m��|�x�c��T�Qe���,��+> ��ˎ쨾;�.�ʊ�x.G�j�n�i$sxj+*�����P�d���[ =M�P�{��S�}���׽]�Do<����̦�ꍘlODCO?������:�H�Sk�4�Ů�R�PK�Ws�@9Y���Rh���	ɛ|�#6����F�"�ힶ������ �r�="��N�)j�4���X�7$"�)�L���B�@����{?ks�E+w��40�`�r��Li�����{�C�ڄ�\�u�y�S?~;��l|nۏu=St�%���Q�Wq��C4�L�MN5� p�Ҳ�h��~]@��X��zƟV�Q��(����ʭ��ߔ�`ˤ���ʬQ��R����o�����O^�~.�2#����6S
��#�"�f2٩`�2�9�n+�8�Mx����8n?�'X��^j����� �;��4������j�o���lai��k��;����4u>d7�Dmk폀�!� U�c�m\�6�x�s��!���Ȧ?H����-0�w�~�H��1ޫw=�!�b��B;s���؟h�GKiu?�����|�5E0��7�<��np/�A+�8^��f7��z�4��R��<���qm|��G�q%\l��u�ev��n��؆4��˸��C�d��&,[\���Peg�T��,) b�9$[��/}�B'kb�u�g�u�NUQh�6��}� �mŨ�ݦ�8��S��с004�L���=��r�[*IGpB:4�a�������>0�WR�$\�&����z��#;6M]���*�/��Ij�1j�ĀR�P3
��7�p��7?#�-�W�!�s��,��Z�2��J?�D�Lb�tu����Z.P��@p�.�}��t�3�߁��	�����\��1Kr
�?��h"=m�6PQ󝠇�A:�~j$pnϫ���R���;+G<B��H3��>s3|�;q יWj�[?d:h[<�v2��� s&+	@oR����%�VV�E�r]�E��X3��櫻,��j��ɤ(�}7o��1�, ���B̖�?���P-�E�[3�Ȯ�1w����T�!G�O}%D{�pgۀ3���?!�]A��U2!�(����Me�T��5�뛕[� ߱N�'�Jh��N�s�2r�p�X�i�C�>�o:�*{�Xb	z�˯sm2d��8�����V�f���tX� ���h;��X��C�x�(�z�� �M��
�hӞ�����Vv�kY���H�}�$U�N���V��DJ��jpX#��G�ɜh\���Def�J ��t_l>� eA��,fgA=��i����'/q�_�2P��7�f��O��9n"E���й����������S7�Y�WK���z���\�ʗk1�?ߵK	�����.g��[�/���HC���.�
��������ʡC#�D��.}x�p(����N�B��y���}�/>�J�Ii�d ��=\G�3#f꨼�,�)?7t	)Y��T�3�$�=յR?Xea���M�z�D�q�/�ц2^_���oų�����류����D�9�H�s��$��?:4Tz�X����9���vI^�)x������Oݟ[���ʰ���9w�`*"V%�zLk9�{cX���k���G�*�FGK�Z{E�*��+�8~�<��ޜc~ �����ǿv.	���u�?�7�/��y	� �B���/߷��h~�}�u���r�*^�X�OP�N�	�����,5kv��Q�Q�)����IO�$�j�[��p5!�6�O�CX����\�[�R����__o/>�TD7�5���Mqè��|��n�~���w�u�f�s&lH�O�P�h=�N^9K�,�����A����͜�	�X�54md���:�!��T#������;|��
y�3����1)xM���8�	�/8�,����w�S����8Q�Ճ
�m7b��ne��eM(���p�|;�M�'g���$�� ��ˁ�l�^�����'���6Wګ����|%z:�����׫�/���Q�VʊSY��);}~�u?-^�b�������T,���:>��bM�-������!9��}f�����9�� L��h^�y�j�1��:�{�;И���Q|�d�r$�1X�p4zgp�-������ܨI8~��ph�w�s��6|e�mH�Ϝ�~'ҧ���R�#Ս_d�Y���}v�j�g�o 7=*%��=�T4t��kJ�h�6$4�A�A�*�V��[I������������*�j��5�W0���T���I"��ӥ߶�'�=�l����%�]DgXS��Ce<�O���j��v�&y�o'R�l�G�C�r�}|M����67�J@��U�1ށ�gW�0��X�O���0Cj��Ҫ玡�J�33�@���<-F��S�����|���E	}%���8�lu�&���<{��O��73>r�]${���"���	m�(�,�,��T!I�=DA5S��b�)&�$J{#��}�0����� ����<\��gg�S��N����N%d�**�<��oDc{U��9j��{�#�+m���X �
IVz�v����ah��|]���(\O`�Y�?���
ۦ�R~�CY-]M<�0/>���#����^b�.�u0�p睾�Vr�9�gb
T��6�{z�P�G����U�ˡ4������'ȵ��kDk/g��Ԋ�끕�R���ݤE�2���f����0(�� �K���.T��r�l'�8�q��C^ ��܆�!ٲu��}�=Ƣ���h,�ԏզȧVxc��uAK���E� �I}���[n���8�W.o��fx~2q�}���9檴�q����h�I4ȅ����7�� TֽG:ʪ�ׄ��]��7���B�:���"������]^ܹ��18P���7`����>�]Gg!Ü��l�!6��w&��c,�f�G*�?�*�h>TW�I\	�7'ᣗ�CI���4X�r�Tl�=��f�V'4���I=��M�Ę",���$ۃґ��[�^�d��K���{�`���y���Ј���=���1Mp��	��0QD-�����L{k��;�4�w��UA0�a��m��[�q-A:�d0fWB�(�'��3�-H<��P�z�I	�^`��o�~d�a�HGm8�4'�q�[�S:�s+o�}V͛@=�B�Մ���۶��e�w�_�c�? �%�Pۂ���}@������i�c/�Ͱ@Q������F� {��w�_bt♻71R{8B�vL����;��H�o�:�Q��`��7d�O�b���`]��'��rJ��%S)2�|�>�K��;��=��h�GR�0T����1���f]����Q5��5Y+�1��|'��f$��
;��U���e��h��?M�?�UR�|�<K5�1Q�OCn�>��KnL�#�Q7�y�ȁ?�Ԏ��2���Ɠve���V���$�Cq�5b%�NW�X�1�:i��F�R���Ɛ��"���UH��`P�k�ef^fk|�qQ��&���gs�9��X��#b�Z3��X%������k[�m��}�"���~������^4U��46�����zj��
�]Q�������D�ǈD���}�8@���M����S��OѩK,��Ʋ��Bt��v�]��T�ע���f�*Y�jB�S�tS�i��.Z�u8�}�;�]�ՉH�wK�F6Q<�U��)��>=�=���)L�и4�՟ �w�F���<Ep����$�
B1�&����V�������Y�z4g��i�uwi�J�f��|��lH�u�
�Pt�A�~��I[��+-�jX�ť��X�l��ڦ=mt������X�Ɂ����b�R}aϹ�v��y���̝�!y�6�N�-x�`������O�:S���O�>o�ӫ�E�zn?��9x�(����u&����
*��i�U��ƫ�����HVc�=������yZE�Z����s?7~Q�r�o$lo�TWl�Æ���cL\O��;,o_y�n���f�8���C^ޜ/'9��P�W�	�C�����uȶ�I?*|����X�^l H�s��$)+*jBi��̌1������-֠ې���*�Q�oO�\������"neY�Z�@��o������LV�v#xo������$�U��5�2��l�k_�M�U_/5�B�����z`5�Ƅ,I'���V� ^�������K��ź��6�#�Ϥ��4�;3E�T5>t�����Z*�SѪl��H�!ac�*uꈉ�>���$����^���ص�����L�k�J��h=�~���Q#�տϩ1 3�:L�-K=�q�1�sP{G
��Vw�0�
��n�f���Y����\�Q���S�M��x��2h���.�<����ӷG�}�hՑʮ%T�R�,{���Φo��[���c)��	M��`��U`��po��yGc	
������YU\�;��[��`��TZ�q�.Xk��XS�58k���<#V�l���%��٠׷kXW����/�׆�g�jq�����8��&]��:�U�~G�X<o��؅Ҷ�1;�,��ᶤ5g�D�ap�AM'�EP�(e�[ 2��k����:�-� �3xPQ6W]>Y�Z|	X���#[�'8�o��	�&��R�(�X� 6{<_�[�������9�F�J!�	y��P����	O�������Zb��U��|)�ё��ϒA����~�2�h��s�j���!������&C����n�F���8��s�=��ϒ/��J9�=�,�'���n�n��������oF�c�,�������`X%t�rY�S��z5+A�I���?��F[��4oT�'U9oɀ&ȤdW�r+�pN	�Pqw���_�a%�H�V����E>R��ke��F4n�p�~��N�߽�QHT��zN:O@E�-��xE��c^�O�����Ti)<��ba��#���><j0,v�s��qaxI���z�ē�Ḧ́�BKCu������B��-H��pbx6�*@�:�/�n?�K����$�cɕ����qy�+��ؙ��C��RfoV��v��}-�=g��v�12
`�a�4S���y3Ӿ���m���,'��fM����*~�M?"/}N=B�I�۪�oL�yݑ4�i����"�����ǧ�!�N֡z�Ŷ_`�a��}�A���g��=�wq�whR����G��%�k=�x�uw K8�s�D���^ԭ`�W�V�nu}T0�&�a�6��k��_�}�xqU|��b��ط��d�o"�D"P<�w�,�L�o���Qp����k�g�m)/�%�� ^Y7����J� ���]�/kh��Z�	�z/��8��7=MS
x�1#/~U㍐ֆUe�-�&�+�6��Y9�2�}:���V.}��r/JBթ�y�)�>Њ���9�bKy��׷�̊�Ԉ[INc�#�gQ4È��A��c0�,HK�2&S�fZU�k���ض�
���J����)>7~;m��^_�U����	���ȟ�P����7�����r����g&c:����6���ݘ94��N��`K���z|w�IkESJ����,$�*fm��ʴL"�)�`kK�(�����DN3�k��T4�Y����v%��`�*��E�nħ�G�Wn�kl��b1���?~�~���Oa�o9W�#Ei��I?��������/�k��o��O�ĸk'����}��tU���`��X��N'�Px�O#*�����t��tX"�5�ϼ��ӝ��D�Ê��S��?��j�&�S�)r�$�x��s���^���p�hy�܂���T��^�*8�QUNw�s|�y�\	)IP�p�
g��m�]ˢC`!�cN��դf�`m-���x��)U��U��|� ��8���x]������rbU?A�"�ߦ`^ �v]�e��
�2���1 Ӕ�y�X]�_:���ՁK��T�n(�M�+��`;:�MH#���=���&m�M�K�B�������C��?��q0
.���̶�.�;A�����(�|�D�1�^Ro�X�̬���)ma<V��'��I���� ������ε�7��<��zrlJ�$�K�z=��^�����3�&vu�3E>K����X�ӒY;�V�e�g��\�#ȳ��thL͖doQ��"**���@�L[���P)f�l��5�,��5�ް�!�T����Q�} !�75�]����]7/)U����ڵ�4;u#씶��$��b-!�c��JU��Q�7�.�Bb�]²	����~o&��$�
��V�=P3�	1S�('��VҦ׃~#�Z���*��t$��<���ݏ���."���s��1�5j�dۖ|�#��8�m�Ƽvs��}}Yћ���f�(]��u�Mt��-���X��R5�s׼o��b��nH���dٰ|A�����0%S�(�q=��omk"��W �v�^p��	"���_p?M��w(G#E��iq�Ut�<�D�f�SQ��mRt	��ר��7�h�	��g�tjvGP9�_�0u'ҋ�NkރU�d�)H���w�A�Z������E���z���M q��f�[p3��������(o�3*�ROC��wlm�sLp�m-�Y`e�0���_�aO��r��n�h�$/�sW��%%]tK|R�R�"W|< �*������˿[Ѭ�u��e�)AO����"��z��Y,��]�!�D�%����eUpQjT�"�)0�����w?	�m���ioM����}c�fij��Yr�Fvqۄ	��rVP���&BBCYF�3hL�Ơ2�g��Ҁ�V�/�A� mO�c�Q��ծ����6�I�=�,�АҠ'̲?���������P����$�&_)ž�e�F9�yW�u�	/A1�hzҷ�-�x�T���'���O�'>]wK��A�	�-7d6��@���9Z��)�X��5!�Y��%��N�^
E jb5��SE|O�SX�'���@���'S��j��9���u��_e�2	;����i["��,-�s0>��f��`6�(V�jM���ӄ���P�q����m]��	v�K����!���@/�-�h<�݁�\ �8z5'�_�R����\������'t���U��jO��h����s�:��P�z+�|���T^�(_\�)^�4�[J͵% X\G��M_��ȽdsS�.| ��o�>�쀨�y������kXt01*&��^M�|�j��Rq�D����͹4��``K;��(ˡWr�!fT���
�>���F�ƈap�&t9j�Tc}lS�f�T�ӆW��h�T��8K� ���G��� �!��b�Pt?��F��Qn�d���T�6'����M� G =-b<o���� �.$���m��X�Sa����a�mh�C �ʭF�`���Q�,בn�`BG�V�uF����>�f����p�!���5G~L����Fw����p<m3O
*��}�A�@@c��ȥ?ԟ��*���v�����⃪��?{�\C��H��Pٌ]I��Wv[]��� ��?l#>y{u�@�����1!�ԁ9�fq�#��9u���sE;y��k�!�-�}� �6�-s�Ȭ%@�l�6���AtZ��W!�oN���E=��$`�3*�D^|����I��#��sot{_S�R�F������R���W�cP�����z*T:Y����o
SlZ6ԋlj���J��0(�GR�r����H��B��I��r���J����+&o��P�e�D�L�� �z�PGQ�&]�à}����Q;v��V]-efIJ0���T�4��.��3&l�u�f�n��n2��X��映��\���#���C�`��/Ȳ�����]P�G)j~l����4?��~�S���t�G����� 5���(���P6�鳮|��t{#���-��� ���[n���(���=��*D��hs(Qe��z����*��f@,�爉ieGM7C ��ڋґa����u��U��&�s�g��V3lb���KC�9j#-�c�H��ߐ��jp9��Iu�V�	'��/T#�Ƅ�~1�6��s�L�,��0]��Iӎ�[ 庖#�P�j���[�u���'IEH�؊�|�g��]��'�C��&��G�U��f�Ĕ$�@=*��O�޸����F[�5M�!x��ƀ�ʜ>�@\GI��zJ\�O.v��).s�`��)r(^��> b��C�H���_�^�!���{\�RLǼ�P�BS�Gsi;��)�^wf4$e79�ESM�@��E�η��z���b�{����#��Sms�rd5�M���Dp�5]��ȝ���{��`.�OK�Xw�I
��ѥuHi�wY���y
['I��M[�@�k3h[�ލ$(�	+{V֗i�F8`e���%b��0%td���u� ��gF�u�~,ӄȺFP�� c�ƻ��xMPq��|z��-�'�39;]_T�5�y�]^�*AvY�ON.~�NU"��|�n�}�u&xU����zQy����F2�9�~$X?��f�����}#P���Y6K�' .��P=Gb�ʫ��ɜ�lI���ݗ�a�oW�����5�8vً.@�GiC�f�AB���7��s-=���/�G=յl2z4}M9Is"�w�TB�3�x��x��t�X0�ٺ��BCH�{]>�@/:N:�x
�>���!��Q����?�6l����ܒ�.U�)B����ehޅd��a,�P��c�͸��wv����qclP)��b�V�V=x��˶p�/}�:�~��ܾ8�����$�[SP��4���5������?ݦ�@
_�=�MM���6[9��"^���p�ߐo�v���s� o���l���"mN[I+A��}����M�2�Z�ɢ�$m.{vq� �C1�X�->kA·�����=$UX���iK�lp�,�C�c����-輨���Ǘ���%]v��?k��Q$ҡ���I�1!˔#J��D%�.��8l6��,O�5�,$��7'Ix��{b/���dѴ�v�`��^�����w=f�E��@e�?A�%tH�=O�������E-&�#	7��Å��@����W*�Rf���afx�bOU��e*X����ƫ�9�]�3f���[�<��z.{���0��F�crA�C����}���\#�.A��]�Y�2`�'E"f���\�s��a8,�b=�9
��A_���5��I7�q.
��Ş�O��Z�\�_j)�]~p*��&�?o�m� ��]\ۆ��)gC�f��y�p�U�#n�{��[�
6�w}f�Q�I����T�Iu���!J���Z�Zu��Y}�m�%��v-�B�����c�{�����1@j|� ����e��Ӎ-���k�$R��C�VC1J��$� B�R�(7����h.fC�-�5�DZ:�e��請M��$�
��D�Ԕ�rV�E[_w��w-�/X!-��OqrM7z8s��%�����ے����aC��3���\�}�'��1�Q��q��pY漈j��' ��G�5P�r�}C�H̽�,��d	y5�5�u��Y�]��MG�Y��C���	�?���eC��K�����'m~'$��]�U5�\ܘ��YL=V���2�"�e
a�CzT-��`{)�J&T��A�	��mʚә,�o�y�k�6y"�XQ-"a78��NC�2R��й��!@C!��C�=�pU���j� ���U�aH[��c������<�������"��3����C���~�j���r�'З�S���A�c��u�f�6��i(el6��F��1i���l�Ƽ���@�#_�˼�KD~yB_���̆���^
@tXv���=qP��Ge�>��f1Ej�.��>Y����/C���!���Ff�4���;�k�RiҚ�h���<DI�j �Mh`5E�S�%3�l�E�M`��Ic�v5B��y^�)���ê���PQ	�����uN"Q���Gc��)�#�V��"�O�Ϥ`	�Ty�(!�s�g�l��c�= �J�S�38���at4����8]Y}�iV6J��O������,b�o0�����fD�S���w>յ_1�(-)�1l}�ݳ���������u6Ճ�����k��SãsehjF3���fע�B�٪�r=��	|<1��~��0#D�Eޕ�h��1Q���]n��J"#���L���ܛ�?�쀗qO�2�цũ��J�� �^'��U���(�G��gSѼ�B1�R��B���@N��4\�V��`�G`�ǧ���E�L�R.��a�\^���7�%v_j(ͭ�^0�ֱ�e�xl��?�S��	2�ê�e ��eAS�*�Lˀ�gZ�"��2,�F�qX�ͱ��y�W�M�����������4?cnZ�=���9�OS�/�S5������^���R}}
{s|������J:v"N�(�R�YbyGIBA���1D��h�����s$�쌂)��*�o����/�����;�ZC�k�Bq�TR%���>��Ɐ��g�������?��
_�>�}�*��]#�'{RXs�{p�f����%:Ohۤ�RZl�I'�魏r�C�F��WڇƲ�zl2�y\ ��5�bz:o�����e���DYcA�=��[A%	�EG�$i=��Ug����׳p����l+����vKYә���j>4s�dD_\Ꮟ�$�m�Z}Q� =!4=���Վ���3��`�����O��	�Ro��ͬ�_֣�3�_O���ԇ�%��d�Y��>����P���K��z��3җ�͛�t��zj$#��4���Ό7����\E�R A�KRu��hH�gڦiw��x���E@y�j-��[��L�{���{�>�X{�G'<�M�N��Vh�?[D>3.��ιn��)��W�M���@����K�»�;1�W㨅�ϸ��n'*%o���)���~�@��}A=t��"IU4�S���|���p��id����.o؈QTo 5�<�i�	Y��.e�ж+���8���2��A��/2J|��*]�Q��k$b���^8�e(�������@X�^�S�}������7y�ր�m�yg ��A�/ aA�b�O�dڌ<��Bρ��v1�w��4V��<ϒ�Ҝ���c�ڜ��wd-5��;K�NC簋M;��5�6�D�n�  �U$�"h��v��(	��Rp�v���0#�� V�0�&c�<�S���q	����Xaie.Hx��^������!���q����'@�4�ѕ�}l��<���t�G��Ooy��fP<��W�W���� EA��_�9�<Z�������k���r�����I~>�z`�w����%H	2�q�K��1� Q<p_A�6��&���1R�A�.-A�6n]�*�*H]o�Md&b"�Ιy��mN����N���!H$	���jV��O2�B�.�u��vD�&�.��hU�A~�gZ-�8lSe��:H��9G�=��\�"�9��	�(�|�4�Tx�����&bK�*ݒ�r���n2y��e{�Vy��ŲR{s�D�n�[���4�9�{.�.S�a�;��|�s�:{(��k˂m��A�Mt��ո�Tʢ́eS�olă{8S���֣"��"8���_����(��[�� �$�&b�v>K\%h�)�AzU�x8�-P�,�aͬ��\�
C��^K��B�j�{-��VI̔�9�[@��R��	1�~��T C��qo��%	q�U��zE��,,�sPtM��5^	��N�������I���aB�� ���;���M
�	�;�I�xQ��G�ԛ�+˫��ÂT�g�̛(�����+]{��+.^L�%Q�^��Ou(CD)��R�.�����������m����G�wqG^�H��;;�/��MC�D��S%^i>4�u���v����.�%���A7zRv�=��S��p�c��*l^G�Կet�/'��)?E�лV& 9b������bd`�]��1���uS�v�k��z�C'��z<�2{ہ�|�N7c�֎��Ws�Em����6%�9�&/�`�n~�F�7��4ѩ:�Ҟ�.����?�P�{��������	�E���q��9�,Ҍ��X��vh˿�Vu�K2�pe���F�����I{��wv�����P�N#!�a����p�;���n/��X��Ϻ-����\Ts��`�_hf�=����8��A��>����߃��-�C-}����" ���7f�cA|Yl�����3��6������L�xd�n)�T@e�6萋rRx��2�G(�85ڲ.K&b��>Xʂ������ϲ�s�^��iW�	E��{�]���|G��J�t{ũ�[]m�QH "���5�d*W%UA>�Q{:�����e ���Qf�'yns۴�v/r��H}@f���j<�C�p�¥�t��B�Ut��
�Gd� *���ԱhTrf��t7�O#K�ݙ�0�&(`��L��{Ϝ������!��QN8ZqP��"A4d��-{D�C�S0�	�m�s�G���QQ�6��Q�
��$�������h��O� �ౘS���oδ�!�1��p��mY� �#�x��.�$5E�Ῑi��&�Y������������!b2OY�m��F�U@����@(��/L��������8
�Y�:=�����U���(�� �㱌xIg&ua{bD^���룆��0�`o9�¯i��3���o��b��D;��������w���R��(�@���(g����W'ӭ R���x�D0��	�+_�1������'Y� ��Go��졵��my�`cTL9E�V�� ��{ ��`�C��=�)���#��
��g�+s��ά��W!.#KV�tK��c3w,����.7L��d]�s>RLM� �o���~t��%�0*q�������<Ga���x�"�w�TViG�.XV��o.w��!U7�h/]���>IA2Y����W��|�Ԧz��t:��y��b~��o#�w�i��@o���)�BJ�[p��h�Q�Y����x��E).�i�y�����*L��A� ��ܝ��wד���zl���u��g��6��B���sG�c�g��� ��g84!{�J�B@9�S�����6�1���D_�:�З^Y�Ћ�
�Cb;��t8�_|�-��3V���~M3��T��wW��0��kkw{���'�\��%�<���x���RT��$=�^����X��un�N�FF�u�#�tm������%������m�q{�2���o^ƾ;1njb�\Q:� ��=B:�'��MӾz�'?T�#a"���d��`���;h�Lt���]��?^�� �xة'��\��A�`|�4Guq�ɺ��}��܂�@�^����b1qV>H��R�
�cS8�~|ׁ�==���ݟ�ߙ	��J��� ��-�p4Q�Qo� �{
糕�-��#�I�8zN����}���O�0A�K�����J)u_�]��ぢ�TE���������l����8�܂񸇔���ggŴ[~��r_V���,;sB��Y��K���-B�LDc�e���m=sWO[KE%؈�يð���ܠ]2������G<5c;/1���ͭ�h��[�F/���3���리H�i.��
~��7%n����?;c�Q��{�1�7aGw^��J"��r��%\$�LL>i{��c1�uR'+ڀ-~&-��R�� ��Qc�2U���أ���I���Q�������(;�y׻O2��7�N	c�<��S�T���2���Z;�fW2VO�xǏ��/�^���'���?M�7��9�)�T�/���k���x5h�4���>�~s�ཷ�����9e��bY�)>_%T� �-7?��uԽ�qI7 .Vl���s�Ҡ!�r �q��q��G�i6���M�Ȇi���4R��#.�^C'�Hq9:��A\Z���a�v;�^/��%Y��H&R*Pǥ����r�mA\��G����:��A���g�~U�id�CI^�n
M7+8���@^F�iw��d��4���Â����X�>��?o�Ǵ#}�T6�L����P]q�ş�JVi\u���+H�cJ�⓶=L� �_ �0,p���\g�d�Q2U�J��#�X����+;�g9�E�5 ���b�N�F�0�!��Si�Gdߑ������f����#�Z�n*_�?TY�k5�G�k:a������a/��.�z!�0߼Oi�*񖡏[��'��N�=`� �+��Ÿ���ۚTL(%�q��"�����x��9w	r����+m<3G���c��"����-�v���Y�;8w�$������U��'i�\AN.������pv|�L����}��!_X���~4&`����x��1�Z�M�}��ި۲v�d�k�ɼ�K����f��ՄWU�����=_a]�x�,������]����[��8��L�W�Wk|�{,�S.>WmTj|v@z��V����=z���1�3L���YI)�(؂9Yؙqz�fnq�a&� �����S��fm�2K�˳@	���ܗ�����
�vp�H��|cG*9S�4�ø�#Kت��V�#>5Aͩ3;2�a����\��X̳�`#�>��i�e.m���ZfD��?5~�
jy1H��Vs-�sȡc�F0�o�Y�F�@w��t;L+`h�6�/qj�sY(�]�N��׶G	A4Ԃ]DQP�WS:0G������e�䆇�.V����g�5��Ւ���L�>�v�>�h 0nU���\���;Ċ����{�o�rA�0Tqќ!����R���|��8����'&|%�.�;t^Ƥ�N�e��?���[c;+�����
+n�5%s�O(y
��"���[��LAR��F���osF��}<�4z
˗~g�!aJ�7����Cl0g��>F�w�r�S@S�{��%�2b�T`�M��ΓA,�Z�8*�Kn;X��k]��Հ�̺_�'�;��:�L�bZS/o�S��G�ӽU��4���0u3��X	k���;���l�@Kd�Lz� ����-����eD��id�+Wgt�ˏ1�Ĕ��pBp�&�,,ʨ�"�)o�*,�'6�&��
~���F��w-�i©�e�j��m�E	�ˋu���{����)L���@�KՐ�e�z��/.cB��ʊ\]�X��<+��x@F�*M�N:1�a�^Ua"��:�;�Y�va�h�/3�y��J�E�~[��I��b�k��S�E\uC�����^�qc�U2R���h=���E+��%��W:�v̅$~���֦��[��=#nb ��@��s�r��1��ZS�U�@���!�n�.RH.���Rd;��\��,�.��c>���i�錎6����z�&�몬AxEj�Da�)��'7Y0�bMx�ן$N�э�@B
�>�y�E��s���[�=|������op�áO/d��^Q�y繏�~u��׶��c���P~�c���b����cr"eD&o�V����Q)�����p`�z1���>7�}x,��9,��t��m�T-�Q��C?@
�]�����4��l�O�"�Fk�ss��,��g����h��.Y�Bt�}U �u0ː���Y��
7/��Kja�O��x@4�	|_�I 0dIȠ;i_���R,+@V�X?Q���e�s�&������"~�Sjn�,6����E������UI��u��5���B;���ܭ�0�ָ-�ZJ�Z�E� =�g1I��݂
����q��5:# >e�N:(X�����FY�.^�����'zR�=��D�|�X?N/tED��:�Q?60��Br��jrBP�xs=�U�	$�✐{���j��*�z�ɕl�4	�>�$��LX ������U���:�������N��(tO|΅8ޘF!�ǷG�Eՙ��6XQl�8x����T�%�c6�8u�2Cܬz�oo��9�R���f���$���P/��iqē�|�T�6w`/��I��~��0��,��~zG妕P��7m!8��%	�ϵUP���nUh�ጤ��&%�Avb���|�8��"��k�0����B��;T<X����"��Q�ɰe��(���Wq<	����ȡ�w��@� �|$*�%��P���:2j�K��&"����>���֓����s��캌�̊+
v)�rk�z�z�	*8��i�ZCő/�\}B�f� ]sj\m�!2�'&�\�SQ붼讵d ����\��n��������HH -��Oe��î@6��d��ľ+�W�$x�k��'Š�A��kΠ*q�´~�ʍY�Ŵ4�f�38a%�D��RD��X*)�6Nk&iR�X�(=����p/弿�#9�*+F�o)6C�1��.2ՊO�^]��)a�/�Ѳ~BI��Y�geb�2��jS!��뤸~�(~�o��m�?��K��?�n���`�c��ɥe'��X�������ʣ|f�@њ4��lˇ��ZD�e�ھ6�]S�T4)t�1���ѿ��+Q�]�7��\Ց�鴄t� "Yr��,B�v%���Qn����?�d�a4�����E5|����k�0��Y��Vz*B�;�iB�.�SU��[R��nV�z�M�c8�q,"=B���Q-��S���	�/-�%ҿ�,/Z.���1��`JgtW�C��r=D���V�]��$� BS"ۈp>�ξ�M"@W+��W1d�ƺ�����[�_"3Fc����5�����w{0x�����2���P���H��=�u�\|NxG[�*�vo	�:��c�3e~���GI��������~�L���:��[�N�����8��+eճ]�S{�j1#�� �zU|���en���k���љ*��Q״���;-�7�|o�Ċ��H�;��@й���j}�k��L��1��V.��!L�]��ӻ�aq�y���h�5 ���N�}��ү��m��L̔˲��'�"���:P�Bjw,���<�E�al��+��!�Ɵ(��׈`ʡӎD��>QD���N���+\<͵�H&����}C�~���J�Z��P&E���S!��	^�=����7GF��*4�l�}��k���Z��n�6�-_�6��cqLD�^�dD���M\�va�٭kEߠ�ҁ�@��癒���z)�|O�Ӓm�v�B�P�e7{����:YOFI7�P:�ۡ�S￹�9.�crR�O\�@~��&�9φ�5&7{�դ[
ʊnM��C��>�y���*��o,$�t^k��#Q���MSt�srI���s�9�	3T������p�,V'$���.\c��o�K��G�8����Gj�m$�Y���be�˾�X��`U�`#�@�qh�b��?'��p�5+0���]�v�'�wjnј�jb�4Eأ<a�)�ӶQ�yN����=���gkh�! 
��G�і$���4pF��\�'����K�eLD�G����W��x�U[�W^7����P�3�+�L�Qq#�x��HѾ� ۏ}��Y %%Un�Q,(������p��-eɈ�e��H���y�Νl���^�UQ>�1�˪A��'i��#Ci�1Ww|UqI��wؤ�at��v-�ȯ?�ڮA��{�i�+��t�����m��3od N�*��w�;�n�BPOn�̾��1���d�ϱ�q-�7�]x�Pp�<�>K��R�E�`���7�/��W�����:�ݝ{� �Ù����e��f�w��!�.o��؜�3�>L�?�E@�>���:��pr�&D8���X�oXY�� @��BM�E'�ɩ�6_C(݀��߸n*Qd�T��LQ��U�i���0}���<q�Z�)�Li[/G�C���!El��O����b$�-����d��8�)���g�F4�\�-�Z�`;r�n��ӄ%��+T����k�þ=K�'c;��y��2,����j�mP����`�yh�.U�7qYp«��L�[�����(q����:ٍr����0닿�#`q���]��"��ꙫc�RT������bG�r8�cN[8�h��a�7���VU�V�:�d�����u��<�C��ت�A	g�Ⱦ۵�fn|����4S���r�@�v��]bB1!�0�e+w�E�g`���#A�>��?~�f�NF�e4��^N�z:�daް�Sm*�P��$�!��Ѹ,�> ���?VJ05Ꜩh<ʅE}pŲ�I�*�����jw)۟z�\r���|���λ�+�<Z��	ȃ�l`$�
Z�P���D	>L@λ�7���4o�D,A��,��ѴH����#w��]�R���C�M-�3Ȧ�b�pAj��uT���||��y�Dӎ��b���ѽ�!��}�L*K�B�$��	�b1$��] 4j��C�\� U���9<���MK;n�_t�~o�k$�H4��1������Y�x�.��d�[�A��~�V��vp���/f���j�X��p{4fV<�����ÐD#FXq��d�0��T��N�(���c��n�����k�
@pw4X���q2�q1j��)�A�I����(
o����N���=��#c��W�G)	�xߎ����AIr���j�;C^䃕1#ܡ6`��˕c�܃u_��F�
��
�̯��`��
U�னg���may���yҕxM��������7HJk��ω�t��9�~�װ��� ��8�r�Q;�-�~d3����:�_�m���8N���3h�m(����Lƶ\K�D"y����m߭?���J6>%�c�|#@�/�n��<�
-~8��L���z[ZU�:�Ӗ��a	2��\���k,!HB�<�ӌ�<�*s����V��["J�ik��M��VD��gyG���Jp�J��Vb��Ԇ�������gİ��*|�ֵ�^Y�ߐ�J-�e��%��j�~� �(_H ن/n�//�ˮn/t�yD]܏�e�ʧ2�Wڑk��e��=dq�L#G%b���k+^�I�2.U6�pyG��pݐ������'��m��5ۅ���fLR(��N=�f�o9>���d�����5m�>���z�;,G>�!.������ƴd.�W�D�Y����c[��Sḡe��/f}SY���O�7�/<t;����A���Tw^��W ��ܢD��� ]"uSM�g�l�˵��s�[f�M���%4B� mD=���{z���f���=cPZ�X^������+N��K�,h5߃j��s� ��ю�����
k�C�
9p*R�'��b��SMJB�c�m��c5���45P$9��O �*������N$���L17�6������W���%�3{����ˎ6 N�I���D�[mR��1X��\AjJ��&$�������ؙi��p��h���B�����PP�yT~SQ�R$�ldB�h�p���@/�P�{���Ӥ
�)H��:�5u�9�X�.Ư���ꝇ�M�8���/.?2Tq�ڙ�E�\H�'��;�ˬ��k���p�D�q�|֫$��n��f8���a"�T"tf>�#��V �9�8S�z��{g�`ݖ�M5���5	�T�h0���t�k=e���
�6�I��EM��&P�5N���\u�%iB�+� D���a��9u��*���	�|��	��ث�@�Dp���b�Ǩ�Y 3V�m�fcθ��0�,h/�����Mw."��� ���8%�|��z�n<���rG�-�H���g�Ofn��#noZ,4} ��u��O�S,$n��	��e��۩�x���	g���]��.��Q[3��qP�'�[�Ya�p���ˍ��X�$ւ��׋Z�%�2���Aކ�I!��7+�( �B�f���-�Q2v[�6�vP蛓>�ɨ�4ǥ�s��yQI|�'�~Fw���O�̈J��q/���]@ٝ�-IΆ���Rؽ3���D��2�=�{UO$��5�����_� ���j?p��~٤"�R�c��q�q ��{���8H��/d�mTr��=�} �1>qa_��������[�}�"��(v��.V�N#��G�pzq�l�~��H��d���R%�ǥc�w=�a"�,��������f���v�V�!����'�SX��2�/���4DlR�9gd����?Y!� M������G�:W���l����,_'�rj�w
�{eʦ�~v�3P��>�Ye�G�%��H�����Ã+[�u��N�~r]���T�^��!�8L:��.NO�쾵��n�S%cː��wG�$�9tY�p��Ay �W(���a�@��n����r��|�^��ۍP̸�f_��:Eۤ�@�e:�`�owM:� �{cv��f�2��d��$�Dw��W�)*�a5����s����T7��Ҭ �HZ/b^$Q-7�'����kN���ӭ8�vNT*Pq�d|W��x�Ќ:,��
��m���6�هx*���t/��5�0A/��g�.��w�X�a���HPI|m6⶝	�r Q7�<t/���x����l#�_	���F&�k�s����\�����B���S��LM������n��� W��������AP3O�lb�$�A�7{���J���D��E2�B����@��������@]���~�ǯ+��Y5���CHY�ћ��0�"׈D��*8"3��J:;Ut�L� M4W�ޅ���y_�N�X���p��I����M�c@Um_��ԍ�Z�;e}P�ۼ��}�X�.�X�����8�ɡ�� ����,w��[��,W�l{r08�VY�� �ZY�O�N�DY�=���aX'�}�׺�(]�H����z̲����Kj�uoz^�ڋ�VM�s֚�.��_l&�'G��?\>XOt�,��[}��Ì׮��0o<�}!����@ ������D�������fҧ�t�b���]���<�6Ӹ�l�c�_�Yh�a��2C���a��c?%��A�W	e<? ���J5ޗ�����<��k�Sk��^5�hҮ3��d�ƹ��qUic� u�Y���4�"x���k���g�aM�\Q��3_bv��nÕG6}��4�����2E��$��"e��8�6���v�!"�����3��hO������^GS�q��yl��,_B*Y�%����yW#4�{�_<�K�_[�� u���p��e�ʍ��7[�׌�?s>���������y���]���3�:|����`1]S�������&e2���A���.�^9���,��2FA`�G�ONNT�"���U�.�[e��US��(ko�<�A�㧌��٤�!� d����z{J��.s��R�����zuy��=�dz	<��c�x�d
��/�ir`'	�߼ѐz��XS#S2���������\��ZG8l�m��/$ Ჲ���M��+�;�R$vi���r&c�׍y]3��Q�/��n�V�����y|?�M��:d|��v�7��Lc7\s�<}�������ur��.�,�[�k�)�+LQ-�3:9v~��sG��w�#k?�[͌�B���N�t�X�� (>Z��3>��q�Bؒ��*�GT�_�)��JCB��d1��qY�����w������.�q]�J�A(�O��3��.�ऀpg�k�3�=�I�O*�rK�@��;�[��H:��j�G��2Bܭ3���kS>���|.���p���>P�b#N�s�p���V�]�x�&3BjF��/]$���=��@�EW��.4#A_�!��ؖ��T����ԣ�4��sN�P�M�Ow�[MF�SC\�1u�ӄ'�zN߲��T!�`���
���EA�%<��t�[r �}d͟r�#ԝH�[,�x�>)�
["�4P�@O��] v��p���љ�KH1t^8=�b��e$���B�.T��tCAs�TLLз;�Z,�ڝ�qx����9���C�3qVsuV[��dG� b��9�J0��q�fQ_Z(����{9i� ��U}R	aタ���f6:d�z|�o�R-�ŷ��ܒ!���㇘0�t�i�/�%����m�V6��n[<���DZd�X�V�)�~%	���ǰl�R�H2�@V�o�k|�S��m�)<�Ƿ[L��z�3���mT3��X����RY�(�������C����9.~6+��c������o���\`�,���-����#�I��W�,-&��
�����fq���n�;@u]U"Ua?��-��Hxj�aR+=�$�U&�:����g-z3#	�Uw7��Ʌ���3�]"#R��NT^��63~�
�K�a��
*X�U�Ɣ�՝��ϊ��뿵���P
G_��d����]7��9I������?�Xh �(���6a��-3L��������k˗����Q<��G��F�7P���m�(Hy��E��0){���M�S-$�7�����f�� ���U�
�2qm�u�)o���N3�)�H�b$�p;|úh_�zH�<+j\OO���ǀ�#���+h�T���/��3v[t��V�.�l�n�_1���-�g�߇!*�;�e��c��P�g�q��p��(]����*�����1�����_�K�4���Ae��,��l�.k|_�ii�X��l`�$E��+�h��;�!�y���K����s�U��:�$�a���Ǉ��]���d�kk Ń���[YߓW1�7���\kq��)~e^���:>�)�kh��^��8������Rݗ�R늵_*`�(�Oh�ҁu?�ü�m�M=���+L����;�@��D���@��&S]�>�e4;i�tX�ݏ���%�ӛz��x������?��p���y�gÔO~&/9C!h*�-�!�a�3i؊��D��|�z��*��i5���Il��=h�8�Wt��ğe�P>��~?�S�ۡ����м�����([c���U�;I�߈�������}'��oK��Ry�G]L��<dД�I��ѝ�k� ��5hFnu�]M���Jy;�&��9�F���&���l�L)��5$�(�cѡ��rmLDvy �\7OL�m����0U�ű�@��9n/��k5����CY3GՊx�ۏ��x�c�ӆdDR�p���)*F��'�S��B��~b>7�F*��N��KU�T��6�V� �/�d��}��ל#���@�9�GYVD%�Y-��iOǲ��uM+�>�$����(��w/q0��n�3@�_�W�R�b%�&���W���ym���⦯T�����+Y��o]!����w8�׎��uǇ?��P���Ѵ\�!z%����ޛ`i�d�? �z8*�?{�0o4�I;�6A����3�n2�f�sB<��.��1,-�f����P@.��%*�na�B�4���g�ص�^�y�9�+��@��V�+�mI�����"\&�g^�A�0����[[�b�����dE�F����m��{�>��7��(%��qn�We%�+��|�ӎI;���~�_8>�C��YrR-l��H��m��To�P��#����Ol�u�]��	�+�����b�lmu�:�w�L��	eE���
�UOz��9t�ԣ>8G�� �����̨��; (=�^� �?�Ϋ��,�Z���zϳ���<Y�fh�R"�0�P��}�Q��PvRF�`�`�)P0�Z�t/P
���H�`����͹ Ƣ_ #������Q�����(��Ȟ+��$�%Z��!0:�X��Ņs�=�#�g� ���o�H���(G�V�b��A�5ȵU��V���>E�>� �K�3� q�H{ME���g�Y�ژm�~-<��%A4FfwK?�ĸl�@��^�SY"�y7��]�W��z�e\!<l)���88ɤ�(%�?ރ\�W>�?�a�vƯCՆK'�\�������F��56��]-!ƛ�8�JY���]
1�
`VU�N-��Xѯ���Q^L�n��0`ɫ:j�Fu��W�T�p�5�	��_i���?Xh�)J�Uz��R8�MA�tҡ*��p@�:����a�==�̒��yM
��q��r�����Ի�;UӼ2r
�C9�;��}���lfIܦ%g�f�?~E���4��`߉�)��"���[��e[M=Rn�\"��Y����f���mMD�C��z�H��Q�g�I*����z�B�c{����2~�nl����6�V�O����-x
2���<������i�<��������1P�ua���(�4��p%�7�C<=��d����$4K��3�_"�5��I��������aU����,�D����a�k��k�z\_^q1���\i�����J��R�%�0�l~wQ�{d_^�qi��(�h�8!�H��$���/���8��޲�5���8��V<�[�ъ�9��50�̹�Cm��o{����5�)-����8��sl�ˣ�E�zt껍��zYP����.��Hv>���z#m~������LD Pn�EI��E����Y$�����rz�8Fn�;֞�*N�K4�g>P�	JbmD<�i�p�C;�2OǀXcW�zuc�P�:SFh�Ѫ�� �ǭ9%�aБ�=��R�ᝳ��3�[	^{���+h3ԻF�o�a�j�~v�5�L]��,|��I	AFTj̦������o�w�b��0��+t<]BS>�Fo�ˁ8��RYXr�o�X�V��ȕ��qZ.~=sQ&��G&�Y7o���,Pf�"�r��̸�%۔��X�"Ul3����x�a�� �������)gN����r��v�R�^&��V֛+6�/S	��	s;�'ZH3���J�g%�B���d����&���n_Pa4PX��������[�Q2�����M�?�I(���Y�G"���b~��h�}����9O;-��䆼��@*��U����mVN�)4��<��w�1`I�g���/d�S4�@x��#B0WA?n׻:M+`'i7��&�םu(���!�F%�|���9 ��@5�k%hP�����fq�ڟ$�����`�ux�M�&T�Qg��=�I�J>v�WBjrT�W�	�~��3���h���p
-��0�Q�(GPQf��_�.dzJ5�����@�󔒉<d5@^Q�*�g�^	��_k'�`��j�XRZb���%b�G��|׮�@�K����_�]@F�=dC�鰂�%���ͻU te��)��_��
��'����I�y��&Y�td�DN=�� ;x�җ�M��O��� ��ͣ���U�D��)y'[wN�ă����L�l'	��3p��������ݰ�~�V'��.���"Ю�-a>�SnAl�[�u>GN({��?��� ۜ44�����3�ܣ����g�Q�!��N�)����,,E�J���tMp�`���q�Jp�8|��e?��e�3. ����,G�Q�ɸܨ��>�pNb��䪜��u�Z��.��s�ŵ�<Q��\�U�� Hi2Z,`ã���u������`�E:<���5:[�W ���u.<� �|z�	�} �V=���
<,��ɬ�!�j,m���nL!v$�~���
�%��q��,�/��%1n�ϋ��,ۻ�}��+�B˗p	���|F���/���+u�
���o�lX*���d�`��P�+�sbPc���x<�@J�+��f�wnd�L�p9y�VʃԹ�\*t�������b�V<^�Q��y�8��~lj��+�㺥=ī��^g�%�O���+����L�����i� �i\]����3YY���f[~��M*ݟR �r~���.�o'Ǿ��}��68��~&
�Ay��L��I�������}�^y�5��[��߂�a760c����7tar��b�$�2�r���:�%����R���� U(~�U���FIP��)ce�q`�0_>a��Uפ*��A,Ĩ�)�����v5����Hg*Ȼ����{�6VH�s���CGh]���~�%ӥ�]8����r���>�t_g���,ć� ��62{��f����_Ѻ���Ţy^�l#j��<��ȚB�Ú�po3���x�6�=���)���ހ$Yƈ2�kA�z���.Y��<8�V�t������9��4cS�Mm�yE���_�iB�e��j�Э�r��eT�J^������w ������Q2�q�r�������p}���|�z�1� �N$ 3ʎ���������'}.ŲƲG|
4W�Om��շD;��>����\�q'q�E�7V�C(#�k����|��˯ߢu��⍼p��C������V(Gw�
_�5�)��݊Y�1���@##Mo�Y���Ɯ�ʧ=���^dP�
W�RX��ea�� ["�-���V�����x�}�s����ی�:R���y�^�����A�{���JU���I|˻`�؎�&��r��T��@�8#z��s%���A���̍*�2�)"{��Q���ɇe�٫�g.��o��W�������w_g�}���`�kBu<z8�3�̳�Q��F7����d`@��2I���)8L�u5{�#�Ɖ��ѡ�0�l��@	R	K=��x��������_��%��9���aG.B"�=�j��Jt��8��x��"a�D�j���k���'G��N��':Vk!h��K�;_�P9n�s1���CϿn§4������O�]({�{�	���B	ރ�j��7����H<�Nަe��/�Y|>��Lr\�$,ۂ9p�K�*���crc�i�D��N�_���wf�����g�a+SE��+��^脋������+���nC(7U��-�J둀4W�c|I���e$�'t�,{ˠˌ�Tam��H��/.�T�`�tY��ym���� �a�JR��rř|��\ͼ?~�oi�1D`�~�!�UE���!vI���0������|���;<����WDH���/�C�>G$�VDP�:�yV��8�鴧�������\'��(�D�
���l  ݭ�5&`1��c:�ɋ��|��<�>���(�Z�c��r�4�Q�)��CYB"��)����LfL�dX���OGw�}(��&��9�@(/Qa�o|�3�_Md��1v3�'3���R@]$�"wB�l�S�1Gz�S[;Q�M�֎|%�*�+WV�w�,5S��)�C2�0���pc\���Wr���pL���e���sd�
 כU#G��|Z�:by8���B&�ݲ��A]�s�RnP�Z��{0_�F��m�C?��������z Ӈ@���w=��RѪF�LV�w3;FU���^I0b"z�*B�]��I����2�W�I.AU ~z�nS�D��,tH~؝��{<A��%E
��L��'�Pv��~��eG��@>`�۞A^mGj�œHș��q��J�!IQN�:�G�#x���+!����놉�D��K$>��!q�Oq����B�J�!�[�lf��ޝ���B>V��KJ���v�;ih�Q������W%�1$	i:0�����f~�,R�Ԭ�#������ِ���r3�'��_��'�~â���=G7��ۡ�T
�eH�ߦMv�ww����WD�p<L�Uͼ3����.��Ch&��|cT�R���?��	��v��I�N�b0� �|}W@�C:>�H3���!�[�"6��[�.w�-a��oRZ{�Ow�AS�����i�7_����)�xX�)E��s�(y�k�o��p�jE%���}/dbi���|\#us�|�U�D�D���7�$T\�Uo�;�D�8����@��`=#�V�ɵ�����@�=6��_�R`֚Fym`��®���T��T�E*LF�s��z���@U��Jc-+m�j��	��'~����t��<$M��l�����N���H?-�&}��~�j�$d���L��y���
A�_�����,��k��lO a��f�9�r�S5�S�bG�/2�z�oJT��=��8\w�\ς��F�N���@�
z�����;i�+�>"Qr$�0H���"�D�[����uEyܥ��J=5��=�U��
�b�f{uw?���x
�d���r��� >�P<Λ�9{Gr�RB�K�R�Q��s��)87/�z,�Q����/�e7�W���]�i�������f_G=@�c��<M)=����6����\��XYY��n1x@���4��5��-|v���L�%��t6�9G X�ջ��O�W���-¢PY��_w��n����H꺐�/C��O.��]<�[Bb�7N&v�v[�%i�p�K�:8-3��^ ���%;�H`c&�
έR؛�}S�2HX���v_��[�GLbI*B�c1�����A�u�sS؞���U���5��;���G�iuP��Ó���q ��v�r���yV���ED,�� �Ó��Zi�f�d�x��e�I�%.�u���]0�.�Z��y���R91��D����n:*�0E`}?�QJ �~c��G�5ALS9ŘF[� ����]����-�R!�?�����}��M�; h/F���f�Kķs����q�f��l}{ށ0%�:�;�J�>o:����;3r���E���
T�p���aЫ��ni�3��6��_�=��p�j�.�1V���i�M8�+���m�{�Ԍ��aXLR�i5���M��	tCM�V+�^LO��u,[2�a������
���RЩ��9�Lm�%	�e��Af���B�Z�@��m�x/��?��2�T �NO����[��$�Ǿ[�V�/&���s2�-�@�!y����k�6U;��~^�S6��1;��ʦ�T);#&2G�:���cY<Ev`�� ���R���_K����s�b��"����I3&�C��U/S٭5�W����4��o,�+Ld�=�{W���k�nN�!�[O�1�{�a�������Z��m�Kxnm��U���Q�װ*r�V0���׍Uj���'�Ȟ���K�
������"h�~l�����!`���]��"�)?�ry.a����&ѩ��L�VY��.9d�����?�+��B͚�ȴ"����X�N�4_[�*�jg|G�}M��q�2SK�����$w��Ќ�e�}�~zm@��YU?
�@���H`;W����F���m���El0y�_�[�F^(�ۑ��X���y����ҿB���al�E��9�({cq����I��T񀓳���j�9ʸT����|�Jf'�s8�6O/�ǯ{�l���2\ `;g ��JК������m��.���Se�B����"/�߉�y���I�r�v/�o��Z�}�e�sYx? ��lpiM��i��A�`h�j��{�}�7�������q��(*P_�b%���F>��T4/���t{��QC�|j�&�w���m��..�#��h��B��/��h5�2{��.�i-���?ɡf���Q���8Rk��ʅ��N�Be��A�o���U9�ϺH+[�_" 6kᴑ:M�'�W�EE {���P�T��R�0����1�ĊDTl��P63Zˌ4X��[�(��� M&�����~=�]m1D����e!�.8�H�"W&�Q��c�#���r�����4���/Q.K���r'���4����1�R}r�U�C�K�RX:[#>�
��H�UF�Xf��}|�IX�uT�mvt_���6NZ>�F�e4�Z >��H w;O˯�I�ٷ��lǃ�r���>J>�ּ�a,t�x���n}x:G5�� �Bwj&����,d�ǫV9j�Mί/}���Q87
�������x[�X�[X�U ��!$��������9q��l����PS$�t,�?
���elƇ��:�<��m5��ms�J}������t�U4��Q�I�d�%u�͗K��T@�E$��z���p�4Z��JКC�j����|#���(%a����C6���� ~/�} z����C��)oU� z6]r�<q/��0 ��e��n��iE��̴���+#tΈ?�x5�XNzF��W� U)Q�a�+S��AN�d���Fܡ�)��O�y��0*NU%F+����r��7g���=���K�7F1s��T/0���P�hd�i�����5�
�Qعi[��q�d��Alq���γ�tŏ��6J��"l�gN��j
$�Zle��Hk;u�Bљ���=:
	3��y-��t�1x����=��YF�|U>�7l?g�7@�3��K����f �
���f�`J��v�1Cd�_#=��WAm�YVe��FKOu������������Յ#$��S����*����)b�z�~�b�vy��\�v�0_� �����3Pm�K�X�.謕SF���ҚKk���
J���:!���#��"7�1ŀ�k3��C!�����b͊q��]������E?��3>�e�xmL!jFEZ�F�+���/D?@�cy�e���ߗ�w%����EA^tҟX�;�u���*�W+����z9U��Ks�Z��`f��%c�>-�,]���6ڧ� q7�	����=�l
�t���51B���q�&U�ʝ�e2�����S�=�6*p�ռ^�	1L�������qX�N�%��X�������o���AA_�J��GV���eAW����2�iV�Z9G�k����\�L�H2,�2���g��+��s���>�D��Ξ��&��.�B�5�8�c�R�w�r��?jU��a>��j���#vZӅqU�in��������͎�R$�	(^08!ɰa���c�xK�taJ"%?6B�je0��+�ӇL6w6�T�����(FD�ɲF�3��s+���v�������MB'��l�e�Ǆi�J����-9Q$_oI�=�`w��^������C%������0�2n�(�<h�X��P�ִ�W��������S {iu��7���3訾&��ԧP�u��=m��h)ڶ6h��J�Ӳ��>�C�&A���g'- B��"`��W!�;�g�cԭ�?CR�Otڀ\�G@�@�8Ka�hh�|�=�Z���:ͽ;�F�yv��H��F����H�;�;)z��z\xY�cG�Ѿ%�cLm"��3ǹ���c�y���GɆ���T8w�" �u6�����?-0m5���"%�|�؜	Ed�l���c+;��0�q
!�7�<غV#�T&��2�4�w��*N�}��z\��t�sn]�>a�׃���.+"Rt�(�lz�o��$���C�r�����������v�v/cWo��886�I�Δ�S&}�}"~��f��˚���oz��TP�s'�jXzT'm7#M�\UV0V�J�<�"��#!d��Dy!m���7�l��/I���ջ��-�D��;�������j�sEg#M�!����amgՏ,����G����(M��	!�(߫�����$uT0�73�QNq�]��0���^"����q���m�E�1�{S��R�Ȏ~V�b����x�Y�&�~��+
Ҋ� �Zq�$\?���l������((]�ۿ�۪3��7��aU����F�P�	Ð�V�>���ֹm�j)����xa��6��2���6Ѥ؄^Z ���bc�᪙��>}�T:KT�j���y�}�&�����r~]��.�	��4D�����Y���,j>�s���$���`@�oq��+��9��.On�[`�� ���q�W'���{�8�Ȼ�%��������WZ��,Ϙ.�vnJ��/]���~3P(`�`k^=���Tz���!�%d`C��:�$LY�0}��k��i���v|�i���R�D���cfQ����b6/s�� �0I%Y(����_6Z]Qg)$�vI�g�yN��D �æP��h�#����3��zC���L��S�F������=�z9�'�W�?m�L�)r+J�V�6�|� {8���>_�\���i�U8ؐ�'�:Sd�����º��hCT���1��k�H�����4D������@���LH���ny�B�h=��
��aRt�w�m�[�-���\��:��p�dZ0)gU�<������U�BU7�U�R���s-a�N��J����6W��V̲Ӷ��B/(<�����V�D��(�Twr݂~����g�M���W���NoI�P����B�B0�����1���oh�s����,f��������g�d]�[r�0��y�r5]%7�G���)��BJك$�= Y&..��+�^
U?Ѭ����]s]�a�ޭԔz��u���z���I���9��kh���]�ߒv��Th�֖
}^��u}���%����v��;V�����о�kC�^���W�V۹����B7�:������ld�2$���<g�zu�*qp��4����������������k�i�0��y;�:��]2`�1����,�|<�س.`���Y�;��Ĩ���\��gg���N���D���{�P%�΄Lj�{1E�!	�h���y�ϩ!���Z�����Ҏ�Y�W2��7�F��,��(^��uЌ?����Qm�J���:���w���Kj�\�2�z*_K㰂yۯ�<�Ol�q�����}(�F.Ͱ9\�C�$�f�te�Im��ڭ	;�v@�f�n�>�������h�+����)�¾<�Fͦ+��ͻ�������@c����&xw����Y���p�(%]���B��$�r��� $��T
A8��������/-�n�4~/�������aD@/��8���n��.�:2|�<�YƄ|I����^�s�E�b��Yٖx|�yy�����#9���I1c����T�b�Con�����U���*��Zd?��&X����wۚP ���հf�Q���ȅ�1'�ӫ�A,��8�����[�N+nhA<�;���8�Y����'�rSI:I���*�{H���\J	�E���}E(Q'���}H���Ġ�>�%D5P�= ���h�ʁ�d��s��̭�Z�����qe���c��e��%��/�ƕ�0���J�y���t�ݲ�̕w�kۃ+��a>Y�tp��CB������y�� 9	F-���l\8h!��A��-/;�AaC�\+�c|�Ȅ'e=_����<�Z���#�t�`^��;n=(B��0�l�~�Pd<���a���>F�Y���p[�u 7�@�z�b9�Uz�>4�7��h8�Fs��t��L�#P��v���T���ԯ�{��J��F�{%�f���=Ǟ����a��ă�*�+6p7b��N՘jz��2��w�>�9,#���,�v�FzD�g�
lt�;ܛrO-ȏ�R9��+������ ���8K��ض�Q������_ga.~$M�ؔ��L�A ��j7�>	��[f�Z�����>T]��RRro��}n�Ԥ��|R���FX�����)���U��$U.��������.
�U��k9�67ʈu�e��t�~0�jgfV�<c$=Y�{��V��id�)�ָ/�{�<�������O��:fF����3�ԭƩ��g�,#$�^�^��s|�C4d������Ra���g�jz3���M������n`	<�\Iie3��D��a=���M�g(��Õٯ��̆���VF$��)<Dn�o���d���A%SSƀ�����*2��ǀ���/>�Xp|�#�*�!�h��z�e0��U$��_%X��2�oo2,*��-E��x�!��%�z�Roe?Rc���mK�>��M�}�ŷ0���;��EGԒwNh������O���֬TcI���t�,̝1�<*>�J�K�R>>-�wK� �p�
��h���a�ā֯��ݔ�~$լ]�p�#��,y"{�������-gfAs�|+����ng ��������v,HΨ?~v���T�������-Ǯ��br��D�2�m:��}�3&W����|�\^��U��K5vX��G���bn����YD�j�l��ǥ�@i^Ly*�I�C��b Uɻt$33������K�=�!��W)��9�Pa���v��y��	��4�r͈h�V>+���,���#@��\�snپT5�m>��|`����CJmx �g���i��O�� �����d^�J:�#xֻ�|l�_�kզ��I�+�=}wl/�h��M�;���v���S�{�o�Zr�تUrkdz��ϛ&��:-�9��I!kr��,��D�-�� XW�G�i�ဈ���}�!p	����y=��ۘ�gצ���U*����qjCRC�'��Yr��7�	O�������ً�j�r'D`��V���L������1}:���DG|�������*�ߕ?��|@�}͇�[��>+�LㄏŭY�����nW5�n
�X<�VLx�t��c E����N�2�:y	�v��#S�� _�\ٔ�CU��嶡���A_V?��TT��N��u�pҰ��箚_ʝq*H|c����7�,����-��HՎč�<�_��fE��+��*� n�[�����b�Qg3���`�g� �|6V(���s�ㇺ�r#&�*��|S��-����M�Q�/ �£	�7��v�L𱈎�3:x�����~����H��D�d��MG���7���}sUx�?���G]��䦺�T�:�������!�f�+g����t����T����_��R� e�T軤��+t�j��.�s�W8����) �2ˆ���|���tw�H3��CN�n�8��j�|bRz�D:��f1]�υH0p��s�����H_�!-A~D(���cȠW�d`��"mU���v-�#ʹ��K3��� ��5�)>���􅒥�����6 ���S%�w�� %�J/~�DX�s	
e}�3XF�!�9�ua���å��_<9�%��:�)�����^��*� ˨yN��y���B#��9JE�U*��bHl�	Xhxi�발H:��y��}��&yx��L_�0�^k�)��S�Mq��'���Y�@���׿�1��#k� E���Nz�荲�����2�6Y7��G^���s�Ͳ����g[f����s�7����E��V�K�)�x˵�_g�%뗵/M�۸_^��_)&I�����+�������X���,�
�jc��,9(V�U�&_ؘ�����$�qe���o�/�xn��AX���A�K��9�z۪������R����c����4�1�M�(w�ƻQ �����z$|�fa��\��S��Id�x�Ƴ�,Fչ�^����uq*�S��v$�=-N�8��d�E�.��9iX��u4��a��]�  �-�V�����9�F�r)���4�w��&���U���۱����y���-R�k�j)�
Dռ�a�}&7y��J�\��҈|�;s���{!?bśS��)(W1�=����6�X}l5)�����}^r�i�z4��L�bgǜ��#� �N��Zg�L�]����:2:ߜ�2]\�6�] 4���@n�%=>��Ъ����e#�i9�!ye� ��)x�)�:�� �����&^n�|p����f���Q���ڱ��-b�G�'�O�7���U����l&^e�>���,�"j�(:=i��YM�M�`qm�U]�Q�wOF�$(%���IUS�i�_�ۄ���Y�U�u�d���/��Q��`��Bt�[:J�1O!I��u�\H�g!�yF�[˺�R�='�kgk�E}�j�@j���Fh� q��s9իh+�i���Tx�.�'�ԃ"�����r�L,G����8�,��p��2��&ݹ���s�遖�=���e�U������L�ɕ�;��4�����/y�QT� ^�6��+��.�PW��OUZ��-d@]E�z忕
�QcԼSr�1u��]|F�bJ �:'��dg���TWS��h1�}+z�u}_0ڸ�L��痯̲�g�e5?|�P"� 1Ɨ(W�3�BW��]��J�vڐ"��ǣX���CS�c�"�>����?�}��3ʲ�:%��N+��̗�H�&SC���5p_�'R��G2��(��*=��TB������h�t䈖"x��U�18QE�L�P�ŷ隹M>ޣ��ۜ}���=Q|�$�� ���bO�v�*�25�-,(
mc��MB����L�5���V���'hRy��Y6�gO��YS��h���l珹>XxX~T~�K���`��,0+Y�΍�'�H�j�k���I� K����n*���lwĕ��=&�l�����6X���Z��w���B��� ��9h��cY� >Ռ���t'�@x͕5݈�z0^�EM�6��L1��_�3,��z7�i�B��G{�_30f;��xP�]c\��}f��.�U*��8_r-{Asu9x]�D���uK�σ�L�h��Ӓ;��i<d$�G�]��mc����H��>WC~E0$ʥ�����u����5(�
�٫��~^�{��˽#{u�(�)�D�o���q���P���b�\lLOS|um|��T��I"�_ñ�W�99A���+�Ʃm��M2=L��o.�S��l�]9['UU�Ø�� ��1M��
	7��5T��?�p�ca��k��3,W�]������U����N�_�u�!�.���f6W��O�O@�9��ydaZi�Ma '�7�p*�(�1��d�?���B9�z�,���"��o��L� c�6��i�<ů��taG3� �C2$�'M�'��48N6�J�Z�	������M �i�Q�'��+�W8~�E&��[���(N{r=��g®�Jѹ�$&!\
��z�^�n�ީ��L#j����1g�+;�����W,�Z�@����=G��Kl�M �v�� �a���<{��\Y9���{�!�/k��bxk7����z:=�;x�Vb��f~/*NIO �M������jK�����2�{�)�t�����1�7f�\S9�J�I�z�7�D?�5/���a��+�^i�u̤	�����o���@�6HhX7[�X3yؓ3U9��d�nl��f8~V,��-/
��֡&�\�8e/6�j�ᬚ����d't���9����2b����4�an�|f���]1e�`�~�f=W;#�B�DD��3�K�����8����dgWZ�����
�T�.���7�A[��՜��A���܄&�<��J<��<Wl�����ǅ;�����	x��m����z��yx�Ό����jv���	��F���vU��`ْ����Ӥ	��9�>��#Ӵ�VI���k�9�w"�s'|��!(L�K	T�Ϋ�h�Nr���2 &���>n���fp���짉����gC_ٚT��SH�`
^(:��L�l)"��S
�oٞqqz�s�k��%�[q8�'��,�_i���Ģ8l���/��:�����^s�J�W�Ac��6$ֆ��,��̸�k/�W��}��#��b�4���|�U�z!�{�������'a�c���bV��1:�F�'������q�<p�1n_�����{lvM#��-H�z�vR|�L�EF��l�+�FN�H�m<����Z�T�!�!7�uϾ��S<uS�)s��q~	B�P���^��.惴�IW"t�lw�􂢺>!�1�OI{��;�5��T�m�A�Xx?C�>�J�V��ٷ�!F�#���N���7�m���߀O��cѫssQ�嶯%֧��}D�>�,�Ԃi�u;�/O�]!<j�rU�28Ib��F�E��8�kb���hwi���L��n�~Ug��,�O1�VZ�����~?�$�.�����7�ތ����Q��3�O�Ya�j9�y��SS�<�-Y	nXW���^=�TP:�'?�I��ޗk�L:U*�ᠮg ���x+1b�(d�����<c��O����0�BǸL�:�C%�B	��*@�vњ~�h��b���Ƅ"�/�@�O01_u�S%���i/�d��èşu�����-��E��bv}f��ʅ���:�����w�����%��fA�0�)�ծ� �����OG9j��Oey����'�yә6(Y�EN�/Q�����X�(^>\ $4�l�Q�upMQ��_���MH?y�ʐ�՝�s��;�}����Q�������Q�vhf���q_o�����|�s>B,�ݥ��4e}����"�
G���^��%,��Kf��L6V��j�
x��I��H!ȭ������
�tyIL���e}D���k�QBi��\8j�uل�XA�2F
I�+�-�[�+�<)��?��ʳ6]���~Kwr�dޤ�@H$�S��Zrǿ�:�0͔&���!�v��l�����9r�RT�Wk_Ӷ�cUe�ϗ���Ő)�䮇�,�E��>�H�>�^W�H�X�O�iL�>כt�I�y��c.Nr��������6ll������61I{�X�Lh�? ��}�E����[�����4nFℌH|KOޭa"?��w�D�M�VG3�����åm�6}FCV&V�}��������
�ËU=N}��3Ky<��t75�9p�U�v��흽�g�s]�����$h��~*�Ȋ�C����iN�з���:i��)��ކH[;�����i_����[���T5!��p�T��GApA��x>z���������au�J]P|��Tv�# 0��dWmLn�N4��ٽ���#���Q����"��^͸A���A<:���L��&���]�C��,�^��x���!*���q�3k|`����،m�E�6��G¾���$�"{Puǡ����R��anv�#@�=�.$���k���ׂ8e��7̦���Z�	WX[#ٷgalwWp�e0�;��D��ދMD� v�8 �T��{<��䉾b5cn��*KZ_�G ̀0k?�UFm6XE�p��o#A3��g�_���뎺	3�?��X�.2��h����ˏ`���0��}���]|͝�8��%�/�4thtN���ڠ��rl'X�K���K���Q��7�ۗ��l��h+�~�(�#�����kN��T~�Y&&ֲ�n���i�Y�\�L��^����h�fY,8x���'��=v	*UUa�s%I3�&8����:�����6Ǌ���dB��a{���%�N<h=Eš�	��.�!S��b4Y�If5H�.�}����&��9�`�]�-_@���z��/+�k�D�������1��;�8２���6� z�T�.$j^��v�^�/�]�:���&�w|9_O�!��e|��.�J��l1f�z��4�zH�oUӓ�d���n�V&��	��~=�g�)�%����f��v�P��@��Y�>�g�_��	��KT�$d�5�n���|�� �I�Vbk�a)J��H{c|.Z�r>���"%�m��Y�;ES�R��OZ��NU��YUR��>`Q'�3�&���D áܺm%�� �pc�Hn�)ve3����?���J��ć�����M��.�g_�p��"�أ�:�;������!����z��<mD���uɆ��N%aV��Q��`�Ϭ���T�q&��,�wG5g8D�����;�rm݄>b�~1a����Efzx�X9q2w�ӏV9��_I���l�f�Iw�8d&��	��[�)�6ܛ4�������5�|YV��l9���Y�G���T�9���h�
�e���#@�Z�$l[���q���x���ʝ�?��F��;�1�]����_+���3T[%3;e����BZ$N�쐂���̻�$��#i��v�
D��gg1�HϚ�@�N#��NH����ON�l��$$��o�s�x�;ʛ�#��8`V�#��`E�󤛙�
��Ǫ"F��t��C�i(���=2R�e���o�ó�P&���I�h�ky���|�q�o'wp[�NQ����ka<�8��L�Y���+�AR��@���Y/ ��3���3��8]������G���U��&�d�5���pѰ�Y,����/]O�����T�\v?��1c<�u
O��K�����j�{V�n/�sNܻ��ϣ�b;hL�y��7�VTS�<���KL�>��Ao�3�_���h,sg��zoC�;���{���q�̓h^*�Ӌ]+,-�P<[�jTJcM�i�kQ[)#�.���D��z���(�u���`~ d覹4�7������H�	�#�C+��f8�"�7��䲫����R׌���$�g�Qk��tEO��+� � >6[ؤ���Ӧ�ʡ������M���� ��(I��E�r%��X����}��{6��ޭ�A<�����d�kn��>����.��i��I���i�j��)q1�g�ҏ���U�����e��dQ�'�*���U\""l�=�C3��	ϳÄ���G�	�mo<����T~*�("RJ�:���dc���-D���<p����d�ӨOxM�a�=���E&�L�G�t<SL�AN��py�сj�1���)�g��Ʋ����v0]�#
�%7�Z0�-zf%ְi�/ޯ	>�ft�á����.f�g;k�,$��5��;vL�.{lL�v�&�V�c�>Q�.H�$@U��v���(�T��xj=̃%��	qm_��T��m�fg�Z�6�ڲY^mV��PϢ�҇��$�~ �&�t���i�2�8�0M}/�w�0��쏩WU���H��S>=Lt�'��
�'�0��^�"��ҲW���pQ�,�DK&�W |�&�;��PF���ﺜp�E���h(?2������Ra�M^&��cR]�R<��W�´as��l�7�7��pDG:�*�~�ݴ�l�𗖞���&��k�$"�7(w�S�U#ʵ�Ʃ��5ա*��ભx�J��(,����yFjPԼ�A��篹HC�RC���	TM��qB�<�#�GPl�;U��R{���m�%'D�մO�
r�b��`}kgp_Ċ�2-��P��r*��۹a�АL�9x�iM�3��Os*sh���p��~<��R)H4�2_\��.��r��xc	4�b�3���S ���b#��n�o��FE�oo�[T�
�kp6��vE�97\�,��d�sa[Py�+O��)�g�~���'�5��������l��a����0����������$J/'��[nv���bk�k�b���8��D�%��B����x:۞���|_qp���ۆ�.3M��z��7F�ѡ][�����Ft�	�<��Vj��k��7׸�]H{l�\��J';�	�z�ܼa�[ku6��I�1����W�^T�#K4N=7e��-#[/���\a)�	�x�J>�|c;��Γ�X��J�Y�J0/����߀����(&�,1܊Z	^w�G��F݈B2 ��;��-��̇kWE|�:F�A
s�7����SM�#��6�Eƴ��L&/'�iO�xA��G�Ǵ:����i�g����B�u�TMFzX�3�I�S"�E�d��)�Yn����+�!θha�`�R���~��˶�`�Eb�m�v=����:�ɰ��Y�SL�t:�ol��;�^�sbM�>�]!�aJj9���+�0H���%��`�n	X���Li�K�&���7yak�h;��މ� �b�s�\� FגЎ>ҜfWf �E�j�1dƝ��A<I�	�L���:�'���)��`]�k-C�Dh�s��[r���������Lն�$�S������A��9e��s���;��<�ts��r���?�g�� @�t߲ZV6M8B��$�9J� ��Y�� ���g`|q/HF؃���nZG����⇶=9_���/��;��uoG\���n#1���U�Q8�(~4�?�j��w��iP5XLZ �;��5pb|U�w��^+E�<Ld�5$�$#��\��I�@�_�h<�`�q�sAL����B'��6t� ��ӝBe,�S?a{un�̃�a$�;��hϒ���4�}$Pzv5�d8�"+YvJ(.Q��o�˄�7_t~`�`7��K�A�[.�BDU�7�`���x.
u8L��w�<#��x��iRI���̐������XtfT}���#����I�(�hm�"�!� Ŝ�E=\X�q"���-5R���e�Y�D�
����y! P���X�N���,�Pj0-�Y)�a�\[8~�7�Pڜ�u���}9'�Z��� ���g���U��}6p�cM�1�h�ʡz�A*%511trW a����v�iG���ļ;�"�2v:���q�Ϊ�سB<V�� ��@e���j��A��M��8"��h^�D�Xen��pw��1�:�ݏ����v��MҔϽa���@)���LS�&����Q1��-EY�|�A}�8��$�Hy���B=%*��7���e��\�&�w���u�p��h1;�^V�y�]���զ��h�L��C��FX�/l�kdwo����k�����ي�ܳ�渎a�u�e}V;I[l�X(�1D��%�?�Ш�Rh�P�̏P�P�i��Ԛ��#���	l�9蓊���:ܢXQ���������-���6A�tc9�;�weP[��6랩Ҙ��c�ӭh*���s���!� ZBe���f��2_����B�x�������3��
������Y3�Xf�> l�Ii��Y���1�rUg�� e�(�Wb�qL��5�3��v�����@h��<�S�h���g��Ax&��/��a�Q���b@1�	��f/Ǩ �8����
g^�<���/�����<�5Z�eh9��p#�����>�2;^��#�:�aHQG�]�;[�V�z���b�W�bG �r�l�����8Y�D 	0��ȣ1x.{��쉀L}	KaTfU�2h��2��	��ܗ��I(�u�����z j��aܒ��wߺ�(��~����9 �)#�̌v��x��n�)������th�� �,.�پ��n��?O�H�Mw��|��ն�x����lqz*G�<^��&�T.��_���)G��YR�����Q�����
��iŁ!+n�~ғ?|4[	pd.+�dAz`�S�U/�Kb��ʷ�w$M$�W�&�z���M�&�v�8�P����:͓Ib�Ues��"� ����5u�?y�jʂ�Ro�ijT���O����(]��7�/,yo\�c 1^P*3^�|��p���@�n �k��;I$�kmGn�� �u�@ ��6W�Noo�U��<�,��zD��Az���{{ڔ2�V�*Kݢ�?r��\�� ]�K�����{V�jw�'��}n |�����A�j&�a��զ[�%�A:���n���1�w�hj����ۘ��ߚ8�#ӗ�K���wF��7Be���? �$1z�K�B5�;�"Z�l: 'b��?*���Uŝ�\�+�B��/oG��GM���k-9�|����l$��B�=���h�;9E楳ڂM��dp��ۆ�'S�͂��1h&����̎au_��M�z�������zy���f��G�k����s�	�}��ICC~
�$5�9[ѯ�u"XS��L��쾉�Y�6r�[s$eO靚��r?�m~�~���d����b�9��coGܪ
�܀�
��ek�<��j�Q��,k4��NB�qw�*/:9<����e]�ͤ�R�Y^��:^�G������!��LADMrp�x_t���g�����Ǵ���! %؎��h���\���%�Җ㢆f!]��2쌞E�l ���Wk�g����~�Ju�(��O�� �/�T�^hu�J?9�K��kG���~��/�H�����Sа�N��;ϋW�o,��`Z��`�09)��T��aG~F���A���d/D_j����,f���$����JA	KD�;��N _)�]�����⒴�/(�<Z�?3@�6�j�3��{��I������/�0ݳ�Dr��a�\�-�nA�۳�f�c.RD;�凜�Z�t��2*O2�>(�P<�#e���l�#���wƟ(�a���+Y�Zsvb��O�\��4r$����pg]�r���.F�~=�����R�B�2_���ݬ��;1jC��C�oS�)+�̠��~����ȼd�F��1wr͜�1�SVg�Ѷ\G4�O��+�U�Vb#��7�%4DOO��K
��E.h���������\ǩ��K�5�����������L�P��\��p��M�D�,��+{��d��h<�h�`zI/�]�-
,(WaTe(Rq��i�v�C�� ���>a�i�E�����r� X���8x���� |�+�ؽ�ow^4v���FT��WE��9�� D�9���b˚��sI�;�����߯I�[�5�}��8Wht�����A5S�N�Qw��sI �� �%������!�a�����`o�,c��Ƭ���c���k��M�HE�+0�~񑿯����j�I|:����5}�s�\�>v��a^�{�T�8�b�(����C'M��&��][S��kC�ۍD�WQ+��=y(��R{XG-����FA����8ΝkH��a>�b�OZa6d*�Q����zaW���Ⱥ�ԣ@����,���}y��u�IP8K�@ -��9���߿U���(}��F)ri!�������qP�y�F�6BOrK�`򸓦����M�|1�L�¤΂������k��\�Cxwik?
n�D�dd&xgmO=ye����ݍM���[84�#��}�8rKZn_���q�i�9�]�#�
~<Ob-}^Б���M���n��a���گ5`�Zյ*\���G�d&q��[j��Z�[WhN�8��9YhA3]��P$@-�@�p!L˞^�
��1��MD��	�,���4�#b��Sh�ys���uR����bE���9�צ�[��qW��F�ޥ��FoJ�x�)Wa3&�v�HY�c�C�;����i�
�L2u�c��%S�җoO���ceL8_6l(=�|�����S��:R"��4(Z<�w� ̈́f���e[�}La1�o�K��}2����~�
$wg+�j��9�%���܄�\�ҩ!:A�F������HRܥ��0.�����P܊T��>�o�����F.���p�e� Ѥ���Q��L|�@RF{R�^���q(�����V�ϥ�r1�Js���3q�_bPM� �2�r0�~!�<��A`��E�Xn�kY��x�O\���h���F� ũʗ���s-�i�T�E���jl�
�W��'.��T���$� {⩞B�иMzL�J��/`�4�:d���%}���R0bNϹ���P�j9�\*t�13-y<��� )Er�j8�:\O����47`?��⚠f�����=�a�����ͧ?)$���i�?�����������"m�(x|Vik�ݢ1�wm�j�>�!�曙_����u��hA4m���:��҈�� ЃX��lsI�6�.�����H}`ȯ�;�� W�����p����O�ubE�@6���
�vnk4��E˺Σ=���>��~�~8h&T��i�(��{�!ݼ��&�t_)�ky�F��B���St���q]Ƀ����Ȥ�/z*�M�v��gW?��fgd��f����!�GIpQr
�LX����.i�0q
��:|�ͬ�P�Yb��7�tN=Q?^Gb:���p��+��7E|�1W@�"�C6M��$�8Jj9����������YѨ�+_�VX��a�[j��3k� �w�3*�۲6z�ʋخ+&�)�}(��J���2���<�P�u����SK��[��iR4��Y-ż�M�5%¶0���V��\����L��8��wJ�I�m((!����X����ݰ~�X�v�9SN,HH�QqMX���K��ϓ��M�@�~��X���3t�Wk���Fқ�we�b�F�S��j��,w�����Z��Q���g��R���:����!V\���d�g�]��A��G2e~fwZ�Ys���ؕ\�t>p�Ώ:��1�K�4���!�l�渴+�,��\��Jq�.�@d��wl�L��Q�(��_ ��g�um �v��p�� �	����'x�ћ*��s��?I��#�����Q���˱c�����p��
�������]^s򋓇Z�Ā�6�;�*�@�hzbvg ���c��$��:��Q��{,d{[�4� ����HL��ɪ�&��[U⶟ ш���J��;U��w���h�_���Ȯ��|��-��AKи-���!<���7�[�G���Z�6�C����s+O�]P�� ��uiE��=crN.��N=Eꞩ�e�J�c��Խ�˵=���y�^�F����X��w��f.������\I�|��khMu�ͫ肮��O�r
@N^>�R�~����\S��j9Iȸ�fjs1d_��v���P�^����W[N���N��}�[2���(��JTíD��阗1(I�r�yo�圶���Uʗ���^&�a���\���k�8p����|rhbS&�����-�/���k����\mٓ�����n��Xmn�ұGs��8�Һ'`�r%j��x�W���,0sf��Ś��97�B����nu��C����g���B	�\�
:y�ʿm�w�@�\1Os��Xj�7�lL�ن��l�/����b�	�K��"@�*8q��{#N��?U�rv]M���K��t�|�d?S�8`��^5�+GW�h��Se�s��Z����EN�K�x4�����!��]�՘�Wj\S�Ua�����{m�a�A��&���E��G<�y���O�3_�r�W	{�M�!y��V��b4�cYT��Q���!|>Ӧp�TR휖�C8�@�̇�j ���Y�����M�,��L��%ۣK���}��`���M�+_w�/����8~ݦ�x}�tN��jV�詏/^;�I�#0��;�Z�Fy�d)��)���w/l�2΀���[��,�]���b<n�����ʐVm��9ډ��mnl��Xi�$w+{ ��<�#�U���%@#��0��.X�c�-`g?�3��+���9ػ���%1��Q�9��T~N���My�a.L��A��;� ���fd\FP��F_��#�������9
���@- �h� ����V�Y���hi��
��q%�����6A�e���rX;~��F-���å"(;z&fŉ�Q�^s4�h*�Hq��P���仳�ؑ�{fBr�A�31x�+̂+p��[L����*�~���z�!����6$%��#8�x�3M�{2��7�Vl��o#�O�}X�7��ω8q�?"Nv��G��E?��hd�p3E��Ϣv[�yCǾփY������v<�� MT�vv>#�����:8����7ǽ+��!˨Y����_=,��F6���c���.}_�QzK��rt���'|0�m`5���k��C�E=X~6��p� �)dˑo�8�Ֆ��nؠ�I^��:HA C��@|[w}�"σ|
@֑�Z�+#c���Xc�0vS�NP�7|�픪��v��/Qz�`me��踺͘�[z�	�X����oA6����<F�J��P� ���CU��앩�]� 6��`�nDk oc`8#zݨ�f�@�yK���^���l|Ynx�J�ԍv��8�p��|�lb�%[MM�C�SS2Ը��\��O�81�P���-�7��Zv�s,�]�{4���`�(�Z!���jr��c?�BH2Oe�E����`��7����֑p���������CЊO;�G���-�)���=���Y����~� ����35���f��b��4����E��4��u9���e[��At FM�?�R��E��Lry��$8"���j_�RZ6��]QM�7x�<�2E�l	]��vD�q���#��m7�K����r��芣��&~ �.�g:����j�#���f��9º��Fܬo0��{�J5f*�Grhz�;���ͱt��Zw�q��s�T���iD��\�VV����g���o�v�3-W��,h���ȩ�Y�z�ZZ���G�}�)V��ƹIj�T"�֙`��Ou��Ы��� [�!�q�z�<�hh�yI\C�ߦŷU��e�C��>�c��k���v�]�����BZ/Zaג�ΕC�J��_"4@���4B��p��;Z@.���?��_\@���6���q�G	o���e�(���-�!^+���lV�5�`o�0����i��A^bg<�acRHw�S�̌8��>�/�0%���NY��'(R�-�r��ő��keo��m,�BQ0&.ђћkS��^¯���*%���F���j�S�Z�!����Ś����B(���у��j �E!�s6��v�Y�1�\��&3$x�dײ����<Sk��}�`M&���]�#Ѐ�1oa9<�3��xIj)�i��GP��2�fT�T�J���m)�ڤP�@�#�.��#�ړ���89�����(�{��}3�3��2/�A-IO{��NX�JB����$OƜď����|���<(�[�3��+���e�s���&F�7��<Y2ZLIc^JÍ�v<��~cI���uW�0~��QJ)��+c�7����ʑ�Epcc� qf$�1����ʝq��tDy���-M����\Z������<V�*f8�KJ��Wo�QȠ���D<8�n�]&�e�gJ8@�'��Lu/���T�G����}��Y���d�͌Я���P4X�5ģ��M��5��@���'�b'�fLM��9��\/�c�͜�ֽ�=яnnq��`E��6�m�_�����mn����䢪!�c:�b0f�'d?+qֽ��)1�F;�����	>�(�%J�����!Mx,5V%~�^�]�V��m�|�-�h�����K��؈���5P��a�ğ{��S֮���\G�����(�M=2�Q�� <��}�N��0���V1�&��:�0eV�#A�e'�4q`�n,l���ʁd�5���\"�S������`$�:������/���������U�gt�d\=��M'���U�Fx��W�G���"�y��Q���J�q��XU�� _y])di{R���S�(z>�[��p"E��Ȝ�՝�dn���`�U1�p�܌��G��2):�	��2��.�;}��M32_�=��m��km��{2W2�IT�J����m����g����9���m�����T���@���W�+��lg��Y��N5.�
ǷY㘫��l��f�V�=���־�$Х��˩�Dۃ�2?I�/� LP��r����W����2�:�ۢ���'\h}���C���tm���e!L�5
r�-��;T���z�C���h�BZ?�{<�wcyo`4ܾ�`�eMU��{�v^�뵩μ�'�E���d�㦧AI��&VN'"k�
�i2K,7�o1��]�����q`�YV��;Su^�g{����p����H��z�M���r�*����*ޛ>'=�=�jP�;��]Qȑ
�?cJl�ng	�j���f�}zzu�R�M��F��U)c�H��Zx��[[5E�~
�cH����o�#���|��t�6�?⏀������e��%��}�e��`'}���N�/���@`
�Ůe�kJ�
��<����]����v*�R��#U�����Di�*�U)x}�:�c�9�o�^q[��6��
=������>��<q�5��~XbNϓ����T>N����G��\4�*�@��s���l  -2_�(��n��|ғDS=	G7�2:J�j>�.���7��rBY��M 8���Z'�v����B|�z��?O�`�}�t����W˭^:+>��Z�(3y}�#�bPE{�?��)�D	�
l�㛛P�����R�}� /d���0�Ә��"띛-�V���:#��R �n����L
V#O3�D@C�L�M��-���;0��J:�����̩ℇy!�j���`.��8��i-�,0<�[3ϣ��7
n���3�֛�̨�G'�Ii�C&�n�?<@܄f�<p,.~�eȵ	'r$E[k~ЙkN����4_���f�d�Q��*�����l���˯�]&yf-�����B��pw�w=I�1vr� �Ew�d�v�n���b�	He��@��f1�Q��R��p_��u��SO<�^�p$$��}\ג`]�H6�4_�f��wF�p�w��f#��U��c�s��0�5x!?p�xmR2Q�+c���em�?�����?V�ۖ�J{v��O��Ki���u�l�`ri�--ˉ��r2ĺ�]%�5��T�McN���C9Ė���<E��xpUx�� ��CP�䰂n��e4$�4H�GIͽ�����;~ݩj����o��&�3��Bd[#�?
pݼjc�{�Ė]�X"W��d��65X�A˺"��mE�5��PUaB ?�����ڪB���CC��i,�2Nkg���H㐊q�p탿p�wC�pL�eb�H��H�^���(�/6t�XJ�Re�]��ݲ���P�ܖ\x܋���B6���T
rZ@�f{/��<t��_tPaj�:J�?��Y��1 ��&|�:�
׬�@�n�H����e}��qj:F�?t�>YD�(g� �-�A�u&)�����B��Y�ΎD:؅� ����P�la��ls7	 kYm�1B0&�.��:�: ��������~pCU�sz�B�a�� ��An��剫Ύ ?p����S��E�8
j��Vo8�,,{���ɰ�C�ρ��hi���?2�v���ISd��6?)����7��0'# ͱe�dm��گk������� M�G]�XR�o��b�|�p���ѯ"Q
#�i��Tg��ᇽ�{ou�69g�!�o���6��M��+�tp1�	C�d^�/�M���g�"��{��� `���3q�i��Jy�.!���i,)�Yv��I� ,��a]��cO���c�XHJ�dWC��1�ʎRm�-��p��FŚ��S<%��}R-���P���_'dk{�Rc��ɊW�+�!���A(�э�8/���F�(3���C%S:��4#VÊZ����p�Qw�Ę~[�<M�K�,3��)���Х%�&y� )�C��U_������d'xRvm���O�3�i}�Y�bE|$;X��w�1�b
\�6�h��Hx��2��ͅl� �63�Z:>QJ>�{$�u�յ1Bv �=>B���a1uG���*��E�T0��c.��#��O���zK
E�Q}˂s�#ݯD	c �I4���ݘ�G�5!eK��N[�!o�T�&�gB�{�v��2�n��
��A���M����"�qĝc=ܹ��@�6��N~���]6.!è���(�K�?�`�.�4��f��6�4�S�A�6�UK���/w�E6O����f��.�r^��c֠,���}x�r�n��s�w�`g�SԹrl(aw)/5�xi×��u8J��E+<�/��o������^�x��j
�b\2eVl�L<��J�����U%7:�c�-��������\�G�D\�w
�N���'~�n����c�p��q� ج�ǵ�$�M;7DG�sX���.˗Dz+��l!�;�8��o�����=�i�F�so��z�6�)ȶES��P�&���7���/���~�0oV�bm�z89���y��RN�k��3'��K�)��{U���iÊ����4�|^7��߽��{Q��>U��0ǅ�Wm���Г��ߜ�؂�Y��<)s�Q��d� ���V)�`9�24���9v�"Ǳ������2�Ƒ=��c�� ��8Z����8�7C�:���e�Iه̿Ï,�õ-I��Wt�T
������U*Ϭ�}��r	@�AgI;� �8w�i���_vt$A�|� U���+)�R]Hkh'� <���K7���g��w�b�����n_&�t��o���Ig�w��/�dZ�N�Cg�b>Yp�f�#�|8-l�3��joP���ż�{F���`#R^�Ƣ��X�̆����v�R�+{��)	�B�ҰM��bE�j�fG��O0r�y[Ũ�&^�O�xT�������ZP`jOcO��ĩw��3=Rc��^Vuk #�W�t\#���G�R�^Y-J���a����S6e�P�Q��VJ�o-*r��J�!Β�&A2e�*�s�čD���t�����1���b۵��E�
����q��z��HS��L�e����&x��hݴb:�;�Q�*6ⵈ`�IF�xi/�2��B�<��,���l��^O�@1Ar�=�!��c���46? (�9U��z��s�Ի��R��G���9��ܲ�8E�)A[�i�j��i[,�s�c:6IՊU����P����>�⋔�g���J���l���5����3��l�K6�	N�Ѵ�����Q*�#�_z�_�9t��'&�Gz0�W@D2A�
�x�y'�O���T�a#���TE�S@N� ���T��u��rl�i�xǩ�Z�����(���`;��z�)u�����~���[U��T��0c����^eM�Sխ�dV���k^Ѩ�M�&�p0�+BB�8�����
���Z�P �=��FD��j�!��|�ZB�E`w`w�L��E���O>)���T�܎��5���N%����E���dW����$���)��5NZ,0|��F���s}��Ǥȃ��s}v�(�.�d!y�Jլ�}y������~"��e�B���}���RtP!
S�cDͱ�<F~BsS2���NoUĽ����h8@VLO�{�q�"Lr1��(P]=@~NJ6�.G�˙j��$f`��\�\|�E��@�F�1(����%\��߮m��O� �oV���wIn>Ӿ-D\���
Ť*ۥ6��Е쏝$��(��͉=�_�¼�yaag<�d�^�C�]I'�<�-����Tg�]eA�1d޴F��L��t����A*�
N���UO��?���x�P��A[s�����=P/��!-[Ա��q̃�c�SY�[X���c�<���uOq+�l���4}�8T؈ݝ�L2���r���+�� 'g�kxG
>�#��G�%��x�B�^r��I1���� �l,1�G�"�y�۪�l}���H���a��i��ue���%~�#�si�G[�]ZX	rv�-��x�=�)jJ=J߄��[ܗ�a&<z�W�rc˘>�ʓQs�2l4;v��BEh�3UȎ�~̹i(��4�v�2I+�M���w�CU��D����x{k4� ��� �~�Q0�]�#���֨��g%�I�5�o:�9�>E�(���ϼ�����P��8�����\u�ZћͶ�@�_��m��/��uW~�Ji��K�Nr�ߞé𞙡�q�8^���CSDB���kc�qWb1�esL.b֜Iv�"Qi�1MR-����H�`�[\���=�O����i|�f%)��sI�%7��x]nA�)������Y�[z�qv"	<ӄ���#��^���=3��'ϔ�b�g�j��	� 1i:Cܷ~n\!Ζ���f��lg���!(4�<�c�%�p1a���H���,�?�~ä�C>��#􆿁?��5Ǹ���O6o����DA��](�9 ��BU��d�^_�֒����!��T2g�r��)����<{�w��-�!nL�줜Xj�_Ե�)GEG$e4;���(_�0l��q`$E�00��0�����j��M+��c��M��G�"﹓�����;��޲��v���p2ߘy���@��M��4�ؐ���58�kűB�s�4||I.(P����0Q�s"$�s�������K_d�z&�
�ˮ��d*��/졦P!�Xp��:�_��Nl��c�kl�?u�~	�B_`{�YJ��=�B��$��Y_H܈��Όu���L_:��lx��u#r��ɸm��7q�5{I��I�n���Pi���I5������͒����h�֡����3{�:�S������@>��1kH����eV(i��ë%P��NI���\辙������e!?|��xn<hl��H���_��n����R<� pJ}���Rs�E$P���T[�i��w*���z� �jLK�r���qP�X�f�p9(
����Q@Q�q�ur� �B��@K5�Md#D�J-O���t1n�AOx#��������X7������;v����%?��C`��.�M��P����-W'�$3��Si�SeO�s��ٹt�����ov(:��~ʹ�!�����2�f�_�ޣ��Zh�s�gL��XOPfތ��l�Y��OyR���}Qy�W�Շ��D������8�r�ܳmGB�[�6vt�,��$*%�1�fmƳ�k�RE���
fC�{��K����篑h6԰ӕA-B���6~��)��O�o/��%TM�K
�D�Y��e���g���;���>�t(�ڻIm?�:մP�^9Wps"�����M�!a<|w[%@9�r�Ϛr�,c3�sh��'v��A��˨�b����'	��c]�߳�x+U8�vz����s ȉ�qhEdx��75����oY�W}�8C+�Z�K�L���z5´y�l���Y���۾.[��88 �ƃ��{Yā�z�����ѩT�%�(D� P^ _̒�2p��*�+�pʗamtc��Ie���'ވT&x,	�.SMb������¢(�3ܦI��c��9&�M��|�S�̓�[3O�]�۝�����ٖ�e��i�~��I�0�(X[}U�a'��Ȃ�V�����h)p�5e��_	EA;^���;H�o8b��Pr\��Y���d���Y�YBc���3���wr�:94�1e�>�g��cXg�?0��'���q\ Ț�1�G�f"r,c��U���Q;L- V�]�Ք�X�<�P��{IE '��`-W�!�/W�r�0.��O	�p����
kĢ���-��1�|*�,�K ����FX��s�uhۺ2%�];3��t�� w˽�8#�q�A��e�B��<�j��i1�^�L$�Wma!#r��#��8Ei�2YW�Fa����ϑ��=@�QTP��T`.��C�y��h-��g{�|p��������UkJ����Lk�r�X#��'}3ƟerJ��RU"Ҽ�J��G5D3���ox��E��%E����y��v��֭���yX5�)���!��si^�ZEy,��E<��5`�'THh���R��v������!Fx��k�?b�?;`§^��t�oI��,��� ���J�����#�|ͻ���w��n��E��0�~ ��d�a��o���ӣ�'E�6�Եh�bUk�GA��ޣyW���nX�|�E+�<���2�_��st��檅HC}�yo^�����i9��ҟƵ�k p�G$Bo���+Er/MZ���e�i0z5�d8H=�Rg�:�����6�r�7��A�0��&��9Ӧ�`����߻Ȥ�����	rB��}͎��"�c�q��d ��ߘ0�	U�db&:�pa4�X�*�)%�GTv�du�o݌lV���+�aY1���1+�k��i�BN�_��$hqr�m���j�#�⯹���;0�U;\�����]�� �c|��,ٹr2N�#z{~H�W���9i�?&� �x0{�AcG�yw����,�n�C9n
���/�-~�ƅw���P�v).��rvR�M�D��U�:m�$`+6���R."���e|���Q�Fh<�PJ~��T�.�쪈�Up�Pԗ9�RfHt[�˩^
�t������rCO��i��rǋC���?�5�l��o�/��CF��v�<�i�;rI��0�m����N�^eG���b�_�MU��&ߜ���N"����Wqi�?����}��d�L����$
ᓊ�6l �j���������1oh�]*&JXP��"öU�fyCb�0`�-QD_�V�N

�,�?���Y����u�O��;[ް_,zw�x�]~��Uԣp�	B|�^8�^�A��BG���m�r�2�L�lWK��=�
mjg��L�0�o����;Ū�2�C��w���\R8*�::�z��݀�H`}ʠ�ʃ�f�ܱ?s*�Q���;�I������hyP`��8���6)G8]�XRk�d͓d�|{q�O�dB����A���;0׃c�����q��[�n虽�qx�����]R���;R8�g��B�&���㖮Y��^���^v�ilV�H+�����0E��Lf���ǵVrsC3q�v��z|+���9�r���.��K��܍}���1]��=�@hC]��/�f������x%Őd�W���6�I]�4�l��q�ۢ߀���/#��]�ϳ#���'>|�G+-wc�"� �S�s�9�Х��O�5M�5䱌��ץy�mU��m�O�Xr���	���)P��p�໱4�jP��ǆh�Ŷ��[t�VQ�}_Ys<�����\�j<IeS��b�䎚h���߽ɻ�`h��j�Հ�z|)c�Iߝ��uJ�s���b�9=���F{6����=͌[{fl��977U��պ�|O�P���[���s��~֧�-���P�9^�'�'��nMVe��g==�Y�~��x=�������a8�?��!1C�;�A|�i[Y���g����-��Kۏޤ� N����s�I�*������.J��a%BF9�\T�X\Hb�i�r�`=��;F�$��C�Nޕۙ^=�+�Yݱ�	�DN7�!<�����K��s�ƶf�m��Ǎ�x�����"]7G�qo��R��EM-B�+4�j��h�K��[���|u����D{��k�e������8����o�s�o!�(���
����RpT��?^Vz�3�zDK�x۹NN?v�us���-��\iz�`_]`�@S�m?���ӰN}�tt*��Ѵ�c���y/����i�S��PEԊ��x��|��k�:����#g:t��g�#�Ho�,�%6č�� rrhtxB��_Z�3�=����^�h�]3"�1��u��	����b;��j�bJ���a>�[�F�ق=,�U|�D:zw`4k]n4�C�K�<�t����ȱR�����.4a ��-��0�~@CN��Y���aZ�*�mS���źV@Z��U�_��X�����A|�4=+H����%��Z��h�8r�;��9=Fy���3�4�q� y�d6��8��P��	n�0�����V񏺫�<�a,I���r`�?9g��-��@Josz�w,׍*>��t�^\^%�edړ�����x�_�r��T���������q+��ޚP[��cXK����*��gl��Z4"_j�����l��O��ɜ4�&5�Y��z�	h .J�' �g���pub��&��;A3C���b��^>bAmI^��?:���Qc�|`b�mX�׬^aA�<�?݌N�2�Mx�Ԑ���_�Y@��y? 3�K\����,�R0lIսp6�v���N��_Xح)�⦎ ��`��<c~�a��䪚7��Uyb���ڈ��N@A��\����'h�������?q���_�,=p�9·Vox��l��ض,H��2�p:��K~z���Yj� �nZ���܎�͙�g5�F,⟋��(�9�j<n����$ �4��Ⓞ����cNa �Κj� 6x��L�ۜ���E��@��ޯ{ɈS�(s;8��X�����h+�@�����(�g*^���@ݜCA�9��t�,����(^9E7<�,5�PpI�|?��TLl��?����wy1��BGOnE���m8���'�rƝ0���1S&ǁ�!h쟭��۰�D����{���Y��r�B�"�z�>Y�3Z�Z�2�"��OX04�6�@>ٞ!&M����)!&�b��[� �-Ɨ93OR%�#�2U��$���Hb����Vj>����b`�����i�������.@��Q�U��F���7;H%be�@Y�C����ƺ��&��2��&��%ӍH讬^\���4��u��.����N��>J$����s��/�W D�~_è��h��}V[?�#=�'�XW�*fZ� �������7fU�vdYejԑ�=�4�'\L&��h�84�c��� �o�L��*��g-��9�RVԄ�s�o��B!A�CNϤc�����Y���p�f#~�_��	�?A�Ŧg9r�[��>f*L/yͭ���Ν��}�v.�R&6�n�IJ��uF8��+�zӎ�fw8�������t�_���o#��j���A`�;C飦XCCJ<�	z\	JB=��Ψ�G+��6��*�j,�'F��j:�L6�F�Z{\���\�L]����Z[�`ɇ^��vl�5'�6lGo������6;Y��6@�)~>\cS�pL�Y7W��{��b��Q�����Ywr3�|�B���~n@��i߈��g�5�w&����T
w���ۃR���+U��V9jk��Ɣ�ܾox�A�x3R�N��C��xGOK�6%�!.q�ɵ>�*�5�F7�OҮث��t���OH�J9���P^���*e�W���G��>iF�0�8By��ʮlWN� .��F5Z�;���r�j�8(V�����(1c�	P��ӌt�-�5tA4��A
rgdP7��~�Ӻ�BM�,%��iaV�ƐCZ<*� �������g�~��Rzv)�jaI�rd_k����*�k�t�*��"�=�;��I��}��C����kMӺ��\:�j��'�)�{1�;�
�Gzi��=�h�'E���A,^��2��$ELӥ��X�Ĭ��Sɽ
����~��<��ܕ	�_9��K�x���e(���n�y���YS�d���ȥ�Zms��CJ�PI�H'W�-`L\��~J��~fPg4C��`�][���]D�TA1g�&c���.k�lW-���2�Ù<Q�v=���E���϶cN�e_"�L-G8��k���g��Z*�X��{��S0L�^M	��O+����!�{�-P�'M��5'K@�y)ox%�_��n����/�]�܋���]�Y�-Yi6s�`�$$�584H�,�j�?%���JI�~�/%��+�w�����6�U�	K�2�0�[_��$�#�@xtLQ8X%~_�X�*
]�����^�O�|�NO9P9����ۮ�AWS�X�ȍů�����ʪ�\ĒR�/ X/�)1	E�5;��s��&!�Ce�bjA��`>�8�U�⎱�2=.�Ї}F��a�����\|�6����X,�������c�*���HGȡ|X��T"�P�~�o� *7�,��)t�(�5��_��{��)j���EA��ۿ���=/�x��#�b`iu����5~�c���j,B��Π��'zYgg�����r��K�tQƢ�ݍO�\�ݗ3����n��fL?yo�H��P)�OO��D�Í_:�u�,�w5Lʿ�ɤL��}�	kI������k�4$�
�7V}���ӛ���`GDL`P&Gu5]�k@�"���mP�z��Iu;œ��	�*B�Z���&��:0�;�AW����Rm�i#C+��^�g���V�����#_l�Α`^|=`B�`�]� y�����P�O�@��"7���F�q\�x��b]��e�ռ�8�1��=�]i�3�D+�^�/_��uF��X1F�@�G&<K��L*iL�.��b�Fkpo�'MҜy�@<��H�z� �<�.���f[,�t�۳"�~��*S8��W�X�:�D����T1�bc߲�&~Fs�.S�t�3�#~�k�#�d�$�:7dȈ��Q��V���sI܋H������C����@�L�JEϘr%6�6�m��&��B@`����$)-,Km�DDo�N�~�
@m����
ϷEͦ�e>��c����zz���*O�.u�Q�ѳ��v���vC8���w�-�CT��� �j� �<'6�g��^��{w�w��]���J�[xG046�ї���/]��W�(��d����y��Z��cO��?��k�m��^���=ЏU?HW9��3on
X���M�v�ԡ����RAN폔�˃�6/�~C�Lz����t�]Za���3�\�&�Ꮽ�"K������bj�+(����q�[��Q��t�3�ٲ5r��A�� �>�~c�!�����D����J�Xz6�e]\Pg��-`��	����o]֛��K�34�?U�"$[�m��$���1�.+�F�/�x�ɮ��M8L����$=�Fs�STú��B.���KL�����S�w�b�Ȉ������t2�f���J\pt��/G��-l�$���I���̢ _/ޕ�ԓ۾z�R�D>�gr�/|٩H�s� j���Z��;aĺ��.R�{�{/��t�ۂ�(�Y���g�>W�^�a� 'U��ݒ��g}�^ѵ�~P"B�(Քauz�Jo�K�.i�{o�_D ة�|NcFT�0��|$����JA�@�ŉƆ���=T㜃�bI����v{�)Gf;p���.h=h�=���k�!�Ɏ��:�4�&P�ഭ�E8_��̅�}� �3����"��U������߯Q@<fL�δ*l"Sb����Ƚ���r�II�	lz�WT��Wxi/�94�/M�d���,�,��t�+y��!D��K�}N���#���x�c�MX���y���0�yCl�\)@�G�@�X*F:�ȍ��Z���U��|�
��ĸ@�Odx��2�T��nc �K#�/~�.�ޔ%$k�23 96�����u�HaS��E���l�~�����H�<�<��,�W���}�Py�O>��
}W�u��D1Դ�8��KB�ԩ��}��n���֩�|����^�2�ho���`���6R���f������<ݔ��k D�[$�Fj����3���7o���^AlGTD��	�Bo� ���Z����'+I �=��]�BQ;���p�����b�HO�:��Ǚ5�0����o{@nҟQ@!Bh#L)kR��E�����>�&G�Pp��DD}C��>cۀW̪��8^�i���H ��v�H��6t��V,���������Ί�g�e��c���L���9���|5��J���QP.�>�~���h�/K3Y�ǹU�|�����
y�OO�a�YB
��&�!���_���C��Z[��Eg
u�5Re�KG-g�}<t&���/ݓI ^��DĩR�;.^��z4x1�EʻX�Jj0����fi˘U�~x�*R<��hű�p�m��n�'] B�݉�~�s'�9�F�c�����^��26�=��,�G�5WMӤ�`���"��K���"'B9D��[�m0b^G9s츀�VL��\�;�������ߍ��.�
@���8�O��V�aGޣK�~=�O���ؼ�D[M���0%z	��F�s��Q�#�����6�/:V�J��m?����3�� m�� �J��3¸�w�M�� �/�^�s�w�`FsZ�Q7ch�H�NF�*��s�5[��O�	M�a��e��h_�ف��(^p��W;i��V��}f�M�|�� �S��f�g�1G��^�(z 0d��&H{qu��j��{��$}�bA��|Ǆƣ�Y�}���:�g���:=$b�g��;�I��UI^KzA�!��akړ��[[��Nw\X>6��:R�C�ؿ�n����}��p~`́��v)A@b=v6�W�l�ΒeFНxM�[S`���o�����g�ڮ�]��k�Ca���4L4���Q~���	�+w������4�[
�w�_��8�wr�r߻��F�MX�֦4D�60�:9�E�y��|P���b.!9�k�D����T��[w��>�����g<4�.[|`/��G>�J�gx�r���!J�RY��0�T�,{3�%��m�ɳ1�-������E�:�F&Z����~��T����08t%�{<���݉A6V=���s���}:��(��l@,q-�n�]��w��za��̣����pை�La�e�J�Z���%B���Z��A��m|�&�4R9�3���ZI��9F��#��Y
Pr�����1��:6���F���4d��|�|bGǖ~�����yW�nw�9��4"8�*�~c�Clz��h�kj2����~�+�I� ����íC\n)�?��l�Jf����=�*0��G[�f2�o0��S�jD���䴜lCt~�j�6UBﰸbVeˣ�o�(���ݟ�8��7�<3�0���\﵅F����v\Y�:�Z^�<5��HH�0��!E4Q�SF�йD�VTXi���R^��Dy�#[%݂jbr%��4^v�2Ef�����&���	1�`=+�|P��h�|!��I��*ҳ�����@�[bi��3����De)�/u�	`ې5Tl��%���9� y����� � �f�hż9���~V��gM�M��5��f]��"����h�6�*\wRȰ|"�QG�[2��z+�x�?K��jcl�L�5�|6���� W��3Y�_���hC7���$��bz�2Dp7��|��}�V�n���t�v�}RO��+��&S=��R�Ş��<��z3�t�������u[o�r��Ё�L��*����+�-��F�އK٤�R!�Q�9�o� 7c _$?��d��
0��N��s��"}7�V����%ծ3�OR�KK�����*��2��O'��ɚ�I`?̭�v�o,��Z)�ǡ�ף�i�$�zմ�&��lJ��ґ+Gs��t; ٦7�-����]�]����d����1��~�$v����č!�Gs��!4�|����M*g��/J��8�r���43ʴ.I�Ɛ"����A�,Zh^����g�3E@V��&7�'�$u�ab��P���C��t�F[���������N����yڐ	u,���La�+T�̛ҧJ>e�r�P����ɔ�n�j�GP������$���؎"�x�G�ʘf�g�����;���-�EVN�����{+���o���b�D0�J�C�|;�vBd��[Ӛ�F�7g|Z3�6�y���K/��3��
�h�HR���^�g�S��}o#ӥ���f:w��D�k[��Щ�f���r~��>�Mc\�/�G݉��a��4��g՘A�<�U���F��&`U�"��H��|�Lw0�u,r�L}���2Ia@��KH1���Rf݆��}�9��z���Spc䇲�-����/U�
���q��)#fR&��y�-e�Ê���EL\=੟�c���G�T�,L��\��<�Q�)PZ��W����>�������n3�.:0,'���^��r0�	����CF�viP(�l��â��E�z���}u'Zs�/O��^4R*��Z1gtW�#zi��[S�P�hMP��3���P���R��y����Q��rG]E:�Jv�Q��bGY�����#
��.;Rڧ{�2+�΋���F��v�����?ח�W`�ՙ ���5��b��� @��ȇ@��� :� ���W��+[f�6+^�^)�yX��T�f���@bC�_\�}�]��U߂=g� ���촖*N�3v�����WP��	�6���������U�e4�G5��a��d�� x���!%mCz�ڃɎ�#�w�-f{|tUu���aR�il�L�Q�7"�O2�7�ry��a]�Cfxޜ�1�J��i�Q�N3C��p�89�����X�R�����/�����<��%;�c�dٞ���AhgDj|��5�Sԉq0^A��;p��M��3 �����9�"\꒿Lj�M�oq%J	m����D���j)�B�����:,b������Ua:�Lan���Gk�'
e����q��K�������?[74Yl�bf��%E�r�:4����n��(��L^QrY;5_{�����OPJ�m���*�@����S�e��Ἶ"y0���f���A��&<�uq$�X&3�S�w��׿%�`"\#O��^�v\f蚔���j^����4�{�(vg�����."X$��'�Y�BR��$�sf���4MM4P�S>�B���0i�dx
��o�X������ �6`�먪L�w�W,5�p���(
�
�{�����NC��+��;�sH��7$fTv1�k5�j�ث$��$AU����l�K(D�[2�9��O�ä�-pT-����Oe>	�=8�C:m	�c)<�GI-_kUd*́�yx�Ҝ�1f�u	\7�e�`��#X$J�Cй��>4�������ϑТK4L� 1j��f(]ԩ�,�j�EP���֙n��oL?��1�=�.5���֍���S�Z�í��Mƍ�`�"lY=4����6���hT9l��'Q�P=d �?t��9a���F�LFXs5@�#\ ��4f=1�e.342I���so]��X�@_�z,jU~HM&ӘQ�MMn�J����K��Z߀y��Y���W��������T�)�7�~T� ���=�Q��K
�V<��Xi��"!��|��0��onj3ח�S	j�m�iO{�S*S�y����Z�5N����d���
7���o�;�fl�b��n���Ձ��}�n[�@ykWb�rdh�I�<�Ό��s�):DpL�SO�k�c>�2�htd�F�Nߴ/W&v3�.�؛D��RBUio��k�I�M��ڑI �qꓨ��݈HO�C�u�7���
���&'����}�R��{�_͚��z�~�N�03G���IE��D$�G�Q=��j�)sty�X��  �3T�T�W2�B]�F`��ϒ�~QH��"���@һ�	j�^��<�e3�Ro�)��5؏Y�M�5S`�FY�_�����M��Q���HK�=�"���v#V!A�q%
�ݛKK������	ax���uHe�F�c�l+��"�q�Q��C�y3by�Z�ח
/*�[�12�l��\@�ݸbcR,�-���a_�'�ٻ`ݓ?A�.����f�PM�Q��� �?�I��4����3fC���ϑ�KaA��iQA��w�'�K�w?}�]��x~������4j���Z,����?��j�^=iǱ��$�h��D�}F ��ZH�7�`��.�u�H�P�
�o�"`$E`������oZT�E����pw�o��j����ٹ���-�VS�d��~�6N�-qE%F`��4xʩ�)�wo�H�װ̑M�!�������Q_��Z;��8oX+��D6딪�L6�6�2�ǹ��T��;��5�,Uc�m�%Yii���|����5���.�C�Q������e��nx�z�L�<�}*{E��A5�?8��f�ǋ�al>�P�.j���	��B��:T!��L�� @3+!	>˩�`�<����mp�L��x~~vp
�ZIѾ:��9!>�1ߗ&��hW���P�Sg���d�IY7���xG����S]�0cpW!��-�}��u�D�f&��]^�+���	\z*!A��-��׿���"��!��;��*�4�um�2����L��f�!�����8���<��i��hR���8���۴��
訑��L�{�m�מ�+e�6�oh�0��J�͆���=�c������_%�T�Yv4���%�� =Gw�4K���?D+��9Y�-�fe���������-̅m����E��m�3�z��s���%�ݣq�N�%7�HB�\���bֿ[!�w�]2%WRK=L��lU?c�]�d)���_���kw %V#����v�.�W��h�SoJp�X1R����˶��t�+���z5r�,'n��}	·�e�?�U�0Q����ޱ\��S <=ម�,;�n�.If��3�a见��zJxe}F-,��lv1�o�/�\7&��2R�?��������Qs�� |�;-����	h�Z�K�+�����M���=E��ě�d;��ݮPR(Z�T�'I�+���#vy0c�<�ѡg��7�C��HkEG��8��;1�2��Az�N;�U�Gt�p �A�:�����wt,�l��O�,J�K�g�k��{`}H��u��%����<W�6��x�'0�����������dA��rד^m�~����<po�ҿ�z �[�Q���8�
�y=!�H�p&��<��	͌�0s��3|#2��<��� F=
��L�3�*��Qa�q~?��[�X�.r`�B{�_4ooG��Fg�{%�*���3Kf=�%�zV��{�1��h������.O���l�"Ñ��d��M��q6��'��F�a�� ��]X�ܤ@�{����;����CsG'����y�� ��|"��l?�z�̙�ȅ�M8p��j�����e̺���F�_Qt�:fEN�{n�U;"���4��$|`x,��_�J�_=I�+���(�� 1��N���c�X谀$�w�(x�b\����A���S�@iQ��;����z��n�TEY��<�|�ؑ&&0����d}|n	��d���H*�C��(�p�%�Qb,NZ�Ou��n�gRM�ٓ��ڻm?�|��y�Y��q$_�$�ۮ�o��u�S0ץ����CB�-��eJ	���׳����&I�"%v5�_�j�9}�t�N7���1�B,К�r����� m�� �MT.a>��uG������'��F���6��KfI�=ڑ��[�D-L3\#����	�i��=�!��I�dA���0z�ݻPJC�yoqS�6^���H�(�@��g��j�Զ�$�٫��׊����M[g#;c�Zۛ�ɃF��2�r����f��k�&Iu={����c�v8e�K'����pV{V���	��)�1���b QA~GX{Nf@ª�<��ȝx(�I&�5y�����mϟ;f��J�`3l��O����TbI�&���&�9��l��ۇ"F|��9�K�.��an���T�(�F�Z*\4�A U�v�@����Jwژc�L�v�41� k��%�%�'7�C�O�����ܥYIn1EB��=�&�x�qQp�1�'t��cw
(�E�X�e�䉀|;��_�.��(���S3���.��ǧ۬_�7�xE)xA�Y���8rr8'���S�C��蜴�w�Z�})�v���UX3HB�6�b�W��Z�Ц����3N Ѯئ|I��R�S�s��I+��Ӓ�M����B���@3%83?���f�I���e���D�&�vI�x��26/�'&Z� �A��Ǽ5���%'a�C��������F�L��I�m^����3k��9 �o�=���%���]TH��2iAXS7������,T���WAK�S���r����_��%}c���Q�+�v�d�y�N�E��F���~��W�h6ne8&%S��-�_�.���Wz�F��V�}\?&_��� ��.<�y�2�IPr���^頤P�\�ek��_XXF�#g��6a�_z�ڒ���F[%��b�q�@Y�=�;�O|̻�@;��N^Ҏ!��,�԰��^Qق��f6�+��b�8Ϋ�VN���}X*����W����r\:m�B�E���%h?!^�r�ajO���A!�~δ1	��.X
����ҚM1l�rp�;z5�I)$Vi�����d߫+��.���	e'��x�UҨo��@��5ct�9ﰔ2�x�KVf��=!Aѩ���_y`CbԮ]0X��ߩ$�s�}B��tL��,f;�s�8��8�v�	�sX�����^��ɨ��B�X��7w0����Z�a�b�9h�M�1��ZH�O��',�6��ϸ"������I�����E�8~��z��/�jE����Hv���/3�/ڛ��HX���c+����.��h�ɮ�.'R�F� �2Cl�Vy6�(	����u6gYoG�E9%�R[6���O��|��JV����`4���>N�y�S��цrJ���B�%�4��t7)�6�$&i,���,Iґ�j �\:r��}k�/��Lc�i�;2z`�Zk�&\�J$�H��/D�>�s�#o3����Jת+d��$j*2��pح�ڲ����sP5i�@֐�x� īO/���ƨO�X�q#���K|��m��xm<�v��/8�b���FhaP"�
� ݇��%�ŎR�������Gb|~�L�}�2��6�CN8�,}1�ҭFQ����������xR�`?h)O0?A���Ж<L�#��ykd�)���QN�+�f4��Ok)Z�𘯲�Ƴv������V��?�*�A��W���?+�)E�ǘi�*���	P�i���t"9
�b��U��A�gt�0��D�D�x�Xw�?��8K٭��K�RPc������)�"�M�F��X�#��H�-JX�O^�w-�.^�,CďW��g4ǡ�#��>,h���׏�	ɬ�y6{TH��g����`.%z"��s���9��?^��.X-�9�,Y�!(�2	yV5���!�qX�Ω1��l�s(,O)���j{�5�m K���ޝ����gŹ����]
 �@KIn�7��̾훳z�έxye	���'+�7�%������P��:�U[�Tʷ\���j��ޚ[Ɏ� kP�^��N�A��@���O��S�Wˠ��d�DL��f�?W�Xy[[�a�,�7��v��.l���/I������٣o%jX�AXj�AM��s�W����F�&�k�^�)>�X�@E,���p��p��#f7�s��W�]����G�褘
����_�ƴ��|X�d���
�j2l��>ag�E ���+O[o|
j�����M�'e�F�f:��D���3��a�}�ȕ��&��@8ar�pj�S�Ѡ���
l��9L�2^�;��'q�dJ`	v�YՁEnHvI"h2��e���pJq�E������X80���Z4j�u&X�;Z��3�^nƣ'����#J0�1ܟ�Q��5!��3��h�~�xMd�.@��b͋�I#S��ԩ�z�E�K�Č������>��K�ـŮ�������lK��ο#v�?�xJ���~·���a&��H�\��n�l��!���CeC��S���զΗ�7���--=�>��{��԰!�f��̡_1�k��j�t)n��@�⍟�Hg��%����]k���ۀ)�����l���un�޼�-?��F7�K �:�X+��X�c�+�H��SZ	�:�%:N�oyڧ�%ٌ*�����������^�`^Ԩ��Xy���iy�;%�ț�[7�͕E��my�U����1d���696��z�z�k_L����r��kc�4}dœBl6�qz�ѐ�%��]�����֮��6S+s���	���#]�� �L�I�KQ��\b��w�����|N�ǕT3?�4Qw����"�a���WD�rv~��+Nd/CX�������K��A_����H�o�c���<�������!�i���Q=��7n&>"��mt�Y���ι[�\(�&WJ;;��S˂:�FINH�ˡxͽ�O�cZ[��C���*���:�Fn}�/���C���~k�����R�X"RУ��%@�ۊ��E���w{k���-��N�-ݙ�����Iى_��"���t��2�H;u~��b]5��x<���J�{��s����2��!�~'��R����J5S~b®2����7K�h���r:}���+A�7ʶ=��\5��`1��1=�)sm,�<W�-��z��	̽ ���h�VPĮ�S�|��.x�My��Z��ﯫ��Mg9���v�r4�2?{�f�<��"Ք�r1K���( �і�˘�N��.3D�@�c�����WU�<`h�0��a Gc���I����m����AO�	-͐Q�kH��E�%��>	R���Q~� ,��K�ڶR���_��Y4���C>�,8Y1�q�1#�����˾1���@n�5-D)�L��f]�M#�_`�%S���$�H��)b�:o�5b��v&,��Ez�Ο�?x�`��>��kt�tm��w{��Q�f�}��:�[	�'z�|�j����pSj/WA��Tx���/�G����N���k>a�J�
�]�6x�?bk�cԃ-��>�H;��K�Kl	�s��0,�Q��}�w��w�f�4�;��1����;��^[��D�����CP�?��@����o�B�"<�4���3|�6�J8_�1:��#�e��M�g=iA<��g�����h����g
����u��l�)����x�<W'�F����:�[�q�Ц�;�]��A��i����6o9)�!i��B&�S�(��NL5��� 4�-�u6�J��lߧ���ͲM��jJ4�k�ەV-��M����[�h�ބe�V+f�M��p�8\D.!|c}�_�%l�� �&�U�4���5�!a�s����74,e��"вq�Y�g#��K�d�k�M^��3֫Q�Un��[� �:ֻ赦.����'�����3S��t�9%�dAW��'P���g*|f%�W���� ��F�F�
��>����z�b�[THP�[l�}�N7�B#6�N��8���h@�̺z�6nm�<�L��nX������7�%�ɓ(�����7W2�I�w�i��,>��4����?�эMR�~R"�~y.~&�3:c(V��3�|n�����bB���o�:9կ���$4��7�y��Yx{�՜#S|ɸ���ɮuH�n�y�J�R���-�;`�A��De�%���i��@a�r@���b��m��I⊃��w؂�Iz�X�˙�%�v�d��x=�����q��C��U��8�^Ur}��ECH 0~��dH�F+�.s[�z����/�]�l�+j�sR/�ir�L6���Ƅ�E+u=�-��@3��ِa�|��7T�2���q+9Ƿ�?�8;��J��i b��H�pg �������?4�8R����O(gWO`T֤N�<��~��>Ε�O'�{$�
wň�QU	Pֱ~�u�b.=-*u!�-�2��A4Az��#�����T�|x_p����#��_�p����~)�r��!��B	Ȕ���d�d*U�W����U:֫��)�@�]��ː޳��[�ɘ�/��*@��6L������X%��_��a�Ϛ��Ya��/JE0��ZNS��������)}����x��|��E�e���x�Ժ�oϗ�����������_[�rT؋Mj�Յ��reǗ�4V��"IGd���=^�T6��<�6�<�+���4�;�,ˆ���& ���̒I��kܙ����X,*hH�!��d$g�a,?_����1�7�T�j�h��}�O+���=�#�s��s��=�u1��-e_��s��mY�����SoN�W�(3�	&rkl�0��J�����>�S��5�ȡ��B}{���?Q�"oŦY`([�3p��!
g٣��}����Ȼ��7ޅ�\i+8��G��Qz�(����|�TU?SΌIt���=�)�B:gLa�������O$�'���@�*��(�w�5��o;�� ��B�G��ZC/;B��0�:�u�I�≋.��E:���������r I��Z���T�*�����p�ƹ;��7�P�?�܊H��b9"ta8�ݜ�V>�0��e�Lo�L�ugF�8؊�ݷ����r�:>��S�ED���݆ä�hu�>w�7z2ߏ6�.jDj���z�-`��Z�7�U�F"᭡@�y���\&��	r��۷�N����:�7��U��_4�p�4^�s��R����Μ���V
�+s���u�w:�;��j/�,��᥃��.�>D��Y�抂�<\[���\�!�?����úўU7�J.Dl�Z-���+�a��r�a�߀w�`�����r�����$��X���	�J
�e�ߓQ�cmhX��1<=Z�(.��1݋����,�	һhذp43�mC��L�>����HsyՇz���]�(���2*��\f�����.��T#!N�^���2%d�d�)SkቍT^z�/p2ߩtR�^iD�<������.
�L��\z(Fp�\�"�8�!f�]�����S�(ý���<�[Jx���&4�uK�=mU�L|#�~���O�?��@��v(����G_j��[�y+��$�x<�!3�6���V�����6���8&���p��x�.��&åJ<J�Z��EȨ���mYnA��c��1}m-M�Pf|��3����ӎ���[İ��G�>���Q�o�k4d����O��R���$]�N�>ɼ.���	y��%�< G[����L���G��Ww���������B�fSm���|�iyт[�7��sQ�����.��b��@H�^Ze����%��ߑ��ϕb"�l8[ �Y�(�坍�i��i��
�-0W3���2�:�^��B�f�ݖީ;\�y�x��.N���<��a!�_Q�D���5t��,o�Y�=e0r��P�����#���Aa乍��aƣ��ט��T*�P��҄a4_�'����Aֱ<:�M��?
3lh��/y�Z����B�)�~�j�E:wS�n�	� �mn�� ���E�pBC���Kg�, L?���s㷥��֊0u5�1T[�	,I�m���&H�=�}ڄ	����7�2^fA�ϟ��Z��eAw���g��C�exCk�R��iv���ಫA�@��P}a(�����L��*2�S��ޕ���2����q=\S��ٔ�ڡ��4ڂ�u��꽖d��
��8��Q�В�KmT!K?�L���G���*+N1"
�%�\0�m�q��a��gw� RK[��(���$g��]���b��G��n`�;f�2��w'�둯��4���:��d��ڴ�s�*G�y෤���/�������`�,nSF<I5M+.����9�������Tg"����� ��=.]��*�[U*�5r���)s�&P/� ��ʠ��T�Ci��4��4yV���Fpo����������9�zu��@;�a���<���}��gH`�aeP�fg��	��iO�e ���<�>���Qy�~���pf5�Ea����X��Vd}s�4]A�������#\2��t�i$iî^�;�ֹ���K��1��c8oUy��S�U��1.�KjCtY���?�Qt��._��ug���E�c����? ͦPh��._Wh_��h[�oQ�_��c��!w�`��[��GH�9�~�s?�|��7���#��#Q�������
��r_e`{e-��<4� ����z��`�¹�V����v�e8��Y?>�.����:5���Y��{��q�҄I�2�el nS��hG`6��H�D+d�B�D���	-ĥ�T��pȜ��Eʝ]l��_	��� Ħk�5oJMŝB	n�Hu�H��y�;a>�{:}��6-ҿ�]���jRa�GH����~5�^�!�`�yC��s�Hz�>rvI� ax���3$��Ě���:k��+�C�Z�}�O�/���-Ǎ���c�Q��(���=���,:HrC����M�~[h�Tr�h\ˮ�OR���T�򌇁��P��z���B�'j�4�%yљ.�?D�sayo�R�z�����������+��/}�'�#�v�N�jn��� 3 �<��S������b�\��ŉfYT��Tw�}Ւ��J$�V�p��F�@�ǙzFv�:RT�4ʓ�[(P�B>ԯ/��ٟ��B����$*�?I`F4����{s0T�`�yW>\����Y@���C5y�k���8�I��0�Г@w��'-��7���#�a�`�&J=B�ɳ����Qf��0-��	�>k��S�0+�?�1m��j�H�nG�*�n���Ag����`[MS��ªΰŝ ��},�M
 V��^����]yq�U)\�/1��q�Ĭˤ�v�dE�ԽX�ld���8xUK��P�_b�����Mk��(���c�T�6�g�e�������ȿH�{n��Kq�0���ێ0��p�g֌P�@7��ި与9��?jM�s�T�h,�hf�>�����G��gc��T-��=����Z�/��Ym�hl��7m$���W)8Φ�.��ͧ�Q����1�� ���~�xxA�����R����R��ZfU_������O�Ӳ��h@�
�?#��,��7Y1�6CE������o���[�A��@Arܖ��^�^!��,H�d�4��`����lhu�ⅧU*J��יu�=�z
$Qĺa�-�B���T%1�p��t�n�=g�F��NA��RnX��5n�X���N��w몌��b�AN�T
�i��ѧw��2R�ѧG�}AP��qAF���w
Uw���r�>~���������:g�ׂ;[�6��re-�F��*~�{s>��^���4�
��.c�]����+��F"|?e$ \�])��o�~ (����z�M_�Whfۚ����yr���'Ry�^��!
���P�B<�'Df������j?r���[	X��QA�M*]�h�c�N��1m�7��n�zv�H�j#�O�{2<����1���!�#R	-C�q\�wd�2:�=��72���qG��#�?��.3���H=;䷼5�5�y���XI�2����#��"k�Jf�(�|OuO�i�6���;)'�_�~k����Jc9JшrN��N���=O)���;s���J�}Ւ�N~��&���a��ځ��v�$�'2!�r���v�{y�(zp�.��#��D_�m����kf���(��B�MQ8.�w,��������n��|Lqy���� �*����
)��������:!j�o�D��E�%����fH^9���m4ȥ���E��������'#\�M鞣T���/`�����̿`R� ����Hs��ܦU�[�>���I3_���X(T��_|��Җb6��5A�Ā��٤	��,��G��Z�:�+X=m](F�$*���]����mQ�֭,N���P�δy�>���{�lz��>���v�zǁ*2�ֲ� �^sr:��d�w=Y������<htT�A��#�n �j��J�u�}�8��|�8����Ѧr��d��j��H��H$N����3�$�/�(�!��:�vp�C�_��vc0o�#�z+�֪���%x��{��v���X��3q��ڵ�$�p�5�5��G�����2פ�J�yC��0�B�:�7�B�ٲ���+ۣ������ή��O�{�.7IQ@dS�/��(�S�����M@��Rvn��͉?�%.� �8~v�	=4�7j�AnQ��D��I�y �r`�h�|�M��%C�G6Џ���h�w��=����?5]��6	Tj�h��O�%�ٕmq��o:�v��%b[�7F;`D&˲Q�2��ϊ��D~'ps���J��1VVi����7�5�%�6/��|f�
#hd�7&�<F�3KH�H�B�鴗LPj�;�C:�����­���#@n�/�֝<�Ȩ^�����|�%BS��(ٕ�ɯ�7��-Y(���dc-0a$�� $
!\�%.��f+�Q���3MY=/T���
��i~�i�oZ�O��p i��E�r
���%RA;��*�(H�\h��9�yp��I��c¼" �u�N��MXs���\b��x�mL$%0�x�v���˒���!m+oy�Z3�]^M�ȋ�{g�{�����xp��������5E���R�}'�3����Yڜ��*�=,R*t���<}o��j��T^Ұc�O�7�����Y|�_��t�P��;�6��D�xB�ۢ�SB\2)�5V�{�,����慯���5y���F��O�`wOSt �چ�$;ߕ��ʾ��#�N�W񀓅�2��UKRkAnj��Ɍ�X9�����I�$��G!���J�Yr�MShc�2[�e���R�%��k���x�ʸ�#w?O@cĚ��a���(4�$
!e� �#�`���B"��&QW�����,����B�w��x����y t=wsW�ר-�.*e�N����ˈ�����w�H�ZсN�W��d��[K�L���s#����`Ӥ�pO�h�Dt2/�ޑ������L��y/8UU; )�O-|^�ׯl�2�9=�E"�F�rIPl��.	�E
S�A��Ri6\^;�Թ�6cJ|�O����Ԅ�tg�K��Aa�f�:����R�ל7�u���o��INƃG��Q��9S��A���yo��* (􆈋
8q�s+��H�	V��_K]�XX=�m?F����4��3R�Ѥ�N��'a\#�PNQK��>�{��p跀���DN���]�~�L=������n,{�JDl4��:L�PC;�������㧣�{S,� �F�ґ���w�~)�v��xg���/�5�Ӯ�d���!/�������EA?3p��4�|�'(p�XX����e/�^멾b2��	L��E$:�4H�6�E�����Y��`�~���LT�'�F��G��DbT-�o&�VYô��v���cd�H��=T��7'�Bqz�����|֯FW\��� �$6�|�U�p;�g�g�*Cf��3��� �� 	/�*�Q�{�]�6+pc �8���SËH��n�]��-'��Z���zc1)1(�4�ei`!�6�t�w�p\B,�2p��D�y?%�b���Xu(��JS�+���:ޝʧ�d��O�c���F��?)���$��H
@:��J�#�[�˙r�y`&0�f�Z_	,o�&[]|j<XA4�v�&��:.���)�:O��Cf�v�	����i�d�Kx'�h�,�R�<�6 �3�]����@�В��P�U�%��v����?gܴ5���b�SX�y�׃i�әr'��ƍ�e+�n(X�k3�	<s�̓U�o�Fb�ͥz�e��-j���VUC|�Ke)���c��y�����r�ΊR�Њzlk��Jrv�hm��A��:лO�wP2Fj%�������1��']"`4<�\�*G�}+������`�5��O�y������,z��	X��/u��i��w��ϑl����BP5�ר9W�)��.�h��m��h�>�=���m�6�X�(t��:>H��rU�����+�j�J6�~t��C������8B8�1�ެi0%<[�����x_j�N���==p��^���M��tu�?V�Ǝ&����Q��(qݨX����JZ� ��ta�IKdV�ފuxu��C��7g�b�����Тn'�I_�B|��H��	���^�R���{����0�������`����P	���&s��"<\�����י�gv1��n���x�J0���h����;T�����4`�~�O�+���{;%�qc˅�9Y��E��:��u�O^lr=F��2`d���f�d��t/7�&��8.c|h�yжͽϹ�{�����lkQ��|;�v�콾�ɩ��y����}��E��*�`徧t�n*���(��9���4�!W8y^��j�����pݮ�S�{x�ͺ�Uy����IN7+ä�P�J��"����Gv�4��Hq���j�Y��o��$4�[����L8:�A|�.�kb��%���3s��xB;|?� 5�ر(?J�)�#Pm�'�E��,�%�\��lR~�;PȈp^���ګ��*+ 	"&�h1�l�]tQf��������Rg�s��?�n:��9�Xt} |����i���,�R��^�ew\��W'��2�u�qY�| �xz��8ZWr2�Y��{�vG7%/*���|�`52Ŭ�8���HlҦ<^)���0,�7ԏ���b�d�i�c�����ۓ�w���g�[і�Z�g��.�xi�G]�[�Si�+Z��_��}�vڋ\��]��oԆ&|Ӣ��pBJ�;h�Ex��_E5���P��.�qք�|[�=����meF��@���f&sH�]����{���-X`�����-C�����U�|�aU�k,���(�"4ߚ9ĢePZ9w��d
� ������	�0:(9�* Ƀ�%v/�g�J�2��0\M%�4�Ak2���.�)�@��#���K��#dR�QzM
�:~����� )Yi�m<�JVxN�T@�I�A�`�ۼl�bx"J�tF̽lZ��IJt���Bc?�~� 8�>nu��!���X�]�z�K�v!�W�q��0�Z� O�S� B;|��c;(iC�ƌ~<�?���M�������3���%��s��o?��)q�����fJ ��Uɚ���PԜK�L�U2�s��������{����q��+��[b�����.����P���������=��}	��2�'�ì`VaY�S�	����e���H������y��\^�]�\n�~�>2)<r8kx��P�]*͢>I� kE���s�r���M��J8K��9���
��A���iW�//���s�O���TY�o��%Y�cN5L�4���"�9��|I2Ĺ�v��BUC#t9�r���9N���gǷ�U2�!��̔�Q�����"����SY�����'���je��r`�vn`y>��pS��ν@��E)���#5)��n��3%�;g���C\%��i��(#�L��G�l�NwgL�����w�������|�S�t�zA�Ѳ�[&�q˗���mw|7�.��1����;��o��I��0�� ��j�p)Si��1br�Ge�N�C~�d����w�%��W�8��Ֆ�S_�VmS�����h�K?�a���a��b>�ޘ��><�k�Q��p�_&r?L���zJ+��ڙ8�%��r�4�'��Н�����^gdn��cAW����|����2�V�'��Rsq=�	]T?�Xa�l�՝�����c4���?��� �$�z�V[#��RR"p?4��w�ʑh��<�,���'��H���e0��%�P&�5m��2y����;ލ���
�#텺�)2�9�TZ���r�T�����sk����9l�x֏��W��3fq���W�ݚ�?�h<RX���,�N�/Mm��o�T:h��]�9�� ���Mߐ�\q�`�7=���-V:�n���6;�f�>�V�3*�u"5�yfX�{��}��1Q?��@N� ���ϰ��}O��ʮU��'>��ѻ`剁QiKw9�S�ZRC��R�ɓ�BB�B'f�?��e/>O��@��8������R�ϐ����A}(��������X��*�1ĝO\�)�}2�� ���O_>�a���-sI�M^�|�o���Łn�qP@Y�˞^&�*�ؤ���u��%��j��xs�UT����B��|G��g��:��_�˕v�0�B�kxh��G61>���k�e�h!�f�񻒪:|��b�+s��˖��%ÿ�&?����կh9�ܢ�/����{"P���8q���k�_�O���͗5:Y�9����1����ĮS2�p1�85��%g����0<l\���l��'8�ѩk�z�>��H�N��A�t�XSj�����q��Ǧ4��$�G��Od}��4C��|�ӍmsWI�NT�+�o����%
�M�f�7S��K�"*!��G�Zr3�{hZ�
�,^6Y�	;P�q)Hd�v�Ҟ�]����#�()eo{�}��ş"6F���F�"�(�픫�C�E����<Z;mXx�@��������zDQ�g,�Pg��i�r[�-�$��ݕv�H�>�r�J݈�!N��8�=0]p䀙K�����ʹ���U�JD�/
̼�"�{�MW+j�]o�YǦ�D�$ Mw5�� ?IA�k
�[u_̩"���
�&��[?�E��^���fFB�Q�;3H.�g�Y��_�ԝ)}�]S������B�sK�����[?����G�㻄ą~vJ�N����X�[�d*��Aߩ�%xk�H<r���/hr<�"%��<BD�L.!����Y&pNlBݻ��Q��}�=�7E�
v�֎���M@�����1Y!��6(v ��������)|��!��A�xJ��-����mއ4X��_�% ��i��5M��������"u�ϋuu�0�l"hTN-!t��8*@���(aH�)�;O��q-l �o;�Cˆf�uP'�Rs��<�oŀ�q-�?]�O����	y(ӆ]dz=�ɀP;��]%�!7�,.��	�}(��F~��Xȴ-A�������kI����Vd[�i� � 9� &�r�[�UH�����E^�vxI�� �m�3��bg"d./�uv(I�$�����_����J�[�i?��uP+)��W
x�R�����$�z*�^���L��SCd��5�Mԗ��`��[��u3{��\=�ѻЏߓ����ꉤL��򱝌D�
�N�W˯.i^|�¨m��v��Ѻen�0V�LYYΒ�0y�e�>~���k�>�T#Ie������*�q@iM"1&�:�S�0����nC�$�Jb�ud.]�,q��_�UA�j�t�77wS�]K�Ab���'������_쌂�y'N�cq�������<�!��=�Pڙ��I�(g����0J�O��8��Z�\�>|<	�(�Vz���K0����S��a�Y�H2I=�o��!��F�`NJ��e��#Wc4�w�h�n�X�����>$���a�w�\�.�>ׂ^��B;����Td��=���� d"Q�L��t��ln3ܾ 4t֋zs�-g}���4�9�R E�ɸ��>�e����<�s�^�%��w�g�,B�6�0� �����T�%'�;"`�-_���R�v�Eu%�In�d��U���W4��QG�oV������	�\'ܷ�� �ns �g;d�6VکyO�QW��D��y��x��Zx	TRA�|���?�x ��͖�� KJc �⿮�_ ���O���.;8xؔx���[���Q�<�wXp�f﯁w� �~Y����@�i.p|�J����<�0�DKE-�5�����r���P/	GLmͧ���k������A5�f�~=�50���WQ��ڟ�1�#7���8%6zr����0R�תbn�WQF�!F���Y\U���G���;���0�t�!�.�k#���c���P~�$	�vf��U�Xk,�4�ᖾz���u��;O¡����5�l$�ܱc*U���w�{j*�0�ի�'5aguN�Q2���[��4s/�w慧�}��Rna7�������֛���g�OQoR%%Wl��Vix �N̡o���1B�1�	[�QK��B8�}�l���ڌp��ړCB��}]�Vkk7�G����Z��fSqq��Js��z��ѓB�4�'����p��ۉ���{���}[�қ>�!�^�ҭ�1�gs6J�_]���s'����*_�0;� �`��!5lEc��6!�E�5F�'�5��e ���%};E����ڼU"鲷�S�����t�--�����N��n�����`��)hPV�"�؟zWwH��x�'������o��?�BEuU����9{��ĪfO,l�ݴ�����2��̨�������d���x���S�O�qaNH7Hm���S��˛���[͑��g�hQ��;V�O%�J���Kxwv���8击I*q�������vv[�ѣ��K07�ϏX~I���<W�j/��Y(�4�r��(k+����m	X�Q�y�p�������0L�-�*�[�mU;Ż���T8��"Zaj&�͸���P?��qآ��[�~l���CPnW#�*Tt�'�+!� �+��b$e����Q� ��O�r$=���:8���n�Q�Q�t���#Z�����I6&x��O�m�B-~�~2��*��͚�!A���%�izBp�@�	�u����4w=���z"�>M���+'.�hHߖ�jQj5N�/\��	'����U�ؤ�*�2F�����טf��\P��\�џ9O9�ۄ��_���/J�d线mv�>�P �הŖd��C�Z�ũ[�h,�ʨ�;�x"�7r`;}éGm=�޹��|ӍO��@�
+���>�&�*g7�xN�А�疂I�����L��2�-��  �717���#B�BeP��)�ɔn����7����+@	;X��Q,:�Ǟ��x�z��:I�/~[t|�����aH��v|�,v=�i�˛�;E>Bi��[�X}";�(�6"�_ԛ�&�b4���t]�nB�=��������~��}��ר�"�96�II���ѽ$щ�6�(�5�!sY�!�ԻU+�g�>� ����n{����[����ǹXP*��_�}Nwr��QY�
��Z���{����b9"�d��D|X��$M������1�*� ]�}22���v��T+��p�h��G���j7��l���@�`$�{����xG`�)��k�	))'L���Ԙ?Z���;
�E�b��� �b0tl�\{������eN:-ݺ)zf;������p�=T�E��2S���%�T�$�^0|���R]�\�X���Dc<�"����Bê1����By5�|jð��J�8�"�6o����4�a/3 ��}�����b�&��Lf��0l}�I�s�k�`�o��|�л4����>���<��o�Jr<�N�B�}��	��%��"�d�h9~5��������Y5�yC��b�G|x��o�%J����p0̃��=�r�]����Ʀ��Ew�X��*]h^��?����C���rƷ��u��VU��F�!x�i�F�^�f��K���IlX]-a�-��u����H��Xp�I�M�-��U;^y8C�Saw4��"o��qNp��=�
�8����r5�3$� }�Ч�iM̾���h��u�"�����6���N����~��{��"A��#��vbd�@��?G��p%���Љ����ϵ��U�u�}��,X��@���TQl�:Zp��wH�qNQ ��_>]��<�Q�?(��w.e��.H?j�݋��( �DO�Z�fV�nt5��&�ԭ"�����s+��L��4~�֗_��t+4���*K�kh��G�����$�5�E����:�3h;��ӄe�+c�}�-�X�4wr	>fY�'�q{v!��m��9	n�i�AF+r�m�X�َgǜyF��e��~�d�T�rTy��{c;��-k�yu;ڂ�į���ٝUqLC��x#���%P0/��F(f�,��9d��~���ٓ��`�������lʱUwx,���R뚉��6��l�A�:=S�O�/~�H�u.�(�8�a��%�}Z))W>�C����Ϸ����]����K����.���H���F;ZG�p����=Q��]V�o�-��(����]����V�>	X!�j���C�dg�-�݂@�A��H@1_n�t}�Z���e�B�}x�ıݠ�_F>Yu���JT�)9�K�um�q��f���w����zP�X�V�:�6C��?u�Մ&H���5�[�'��0{܉q��"w���$�/sۺslvEX]�;h��&��M��<O�F���1!64��
�w`q�A8F��>�[[Rey����p��9̟�-�9�ja'�(�.��Y��a�������� l���#��x*Vp�3�`��5k.Hȵ��{6*}Sw�C�V���x9�o�&�����֙�QP�_%�t�$��@�`�=, �x]�iPt��출K��*:��,�p���=&qd�I��Vˑ�U�G�ƕU5�r�4Sp@	�'�T"�S���b���O��Y\"�Կ�}��7'����u�Ƌ�0��$Z�?zd��G��M
R[��I@+�]6�e<L����N���R��甛+?�9x�������C:;_G�"��ב�/ڱ����mK�7~���z�P���O��ո�An���0�o���*	��;�J��v����?��(�wׇ��J֩�}�#
��C��!cU���y��f�8{�m^�-�1K����W��3J����B�莾�3P����VЌfxgZ!�� �[��&Zs@�(�����A\(���<�a��;+�]�!��|	��X��l����D� �:���~����1�a�FsUV��w��v�2<c9�)X��k2'�q3!�����'Q��J��m�()\����~�΂qM�>�H����bx7s��_<��#�������gjkV�)+���"��+�K�E�:�Ey���6?m�T���Ȝ��H坻Z̤�f��V���@0,�Q�<���;�z�f�SC��\���v��b&���Oqv!�~s���얠GL�y[ja9m��a���4�uUL��b�z�*��( ̯8��6��sK��E�=�0�<?A�xQ)[;GW�g�%�^=b�ڌx+X'q_b����T���'����9wg�b�����p��t�o\����u4��N�p53��e�4��R��1�/ǯO�Ĳ�43ObkT���R�{��i~mr6oL.,/i��ùB��{]i�����8Qe3H���y�5u�=8�Z	N��q�Px0CD� ������������u��wH�Q<�x��q��St��4��#�0pa�ՖS�`Ȼ��ߺ\��G��ӒH ���8�fD�����5�rKj�]�#�9�H�/3c��,���V5�w?�r,�cR5暯�^"�M�qmP�̡��Z"�a|~�ꍬ����Qѝ��`a!iǈt(�W�̓?x��
H�3�/��)�R�n�G@d��:�$^+Q�>���§,p�2�m]�&�Z�L�{�rq�Ŧ�;mB[��!��<�%3X��a�A���a�~�O��rǪ8��qI������f��t;q�}%�H�[��L8�"h"I�|I�������A��>Dߏ����wݿ�-5ް 
�X�A�cl���o�}c��=��k��~��+q�۴�)g�P��Sk���#�Ā�i?�Żm��?��o�5���W�Y��+��.1� ��&��k��0y�[�[�*��4�R�]��:�o���QQ���5����u�]��41�����(ug��;������.��;O�wa}<��)u,�j�F4�f������'G=M�'��	Zm��w.�M�x�W��7�0췎�$�Ps^�� ��m�/�Jɮ�%��]� \ۏ��F�e����ݦ�q��k������T�z��qnz'Ek���QL�1�D4��7�������ocV~hsqOYTa�,i��\�@:8�6�eB_}��N�
�q욵2<�z�W� �?�BH\��96�	U�N��-{�\G.ҡ���jё�XT�Ru.b�c3c�4��(0M�[�˱��1P�0������~2d1fX6c����;�,�[�W�J�+��$t$L�+�@�Ü��1���մ4���z�O���,�aP*r6�����ի:��Er�h�#���x���b�T,1����_+��\�<u�V3,�j��>���:�Q�윇V�;�[��Qq�_h�%���a5��Jwe��zd��M��Dh���x�"\7�(*�� u���)�����g�2��f����^{��`HZ)������h,U5��A5�⭃.�ɝ�� '����h�����y�i���xL��"/�#ϹK�|z���b&ץ�{��P��.�l5BEO�#f�l���ʽ���f��AU���d�e�;�7H'=��� ;���kbX��<S�@�����ͦs���]q!��`��B���P���Zc���|�ŉ;���y��^��EQ9�יW_��CC�'@�g�w"�3[��Y�1�����i�1�N�iEC��eY,��H:��.v��ǌ�sf�0tT��~Be�G2^��߫���*���u/�IV7N��u��[M:Я��O�7IWlV!.MR>�D��Z��cg�\�EG�Ze��2�i �^�s_+.��w��t��;������&Z��z�x�#T	��P��DMp�w�A�3+[A������[�J�~Hv�;�t�. ��ˬ%���?5��|�0o�S����.3����xt.����Ը�n��$�.5E�v���6"���t�+#M�99��g��mj��3�y�V �)��ǐG_����&xl�\��~���!|xA'��rmƌÜ�3R��"#����3������\������xz8���i�6��*uj�����������j��_�X���K�u�t�d���ڛ���
�3����0���>���o�������d���jrߌ�j�����"&�B�=�m_w�U�Y+9�4�B<��tj
�0�벘v�v-Sw�y�������i���F����fw²��L|�C+������e��ߙ���-7��<��Y��:W-t�3�����Ӏ����������E�)x_��c�Bd�-������"!�d��sV�(s�s�ީ��7��������v�*�1�SS9?�=�^����^����k\�p)"��_v��;�;;ѩ�"�u)��ʪ�%���/}N/3p�J���tkю&q���Z�&Wc:(��R*�PIg����v�L��G��/�<�g��tr<Kh5U�&mV�*�S�.O3�V[2D�ˎ�/B���ˇ�T�%Z坟+�h 
��(�]��P���a�6r h�q{Pg��)�C�n�O��mFk���loS @\���ɼRAӋ�1�}���ţ��|�Q�2p�Z�������q��(5�܅-��:��%k���'����F�����sz�hh]��X����s�e��bY�B�Y�DF�T��l�E4�lo�]�7�j-=�G6B��|�{��x�$Ӡ�$̏vBJ���v<��|;�W��dX��+�3V���B�u��K��ٽ��)'%�k��T��x�Q��m�����F9~�ډJ��xJ��%�i���Ő	߳�J,��n�,X�AP'�`޼� ���*�>"]�̓�������yrE��@o��MqnIK��M��VB�q7��}�����ml��*���܅��4O)�Ӫ�!�J�r��t$�]t�f���AVI%ڏ������/Ŏz��*�G\�v�͋����4]A4��.��[���X<6�יx�PPߡ�Q��
��ߞ� �D?n��,M���cb�\A�`�yӌ����#�+(V��?�z��L`N�5���$��Ym.�O)ϊר�հ7��s��2g$w��!��ѱ���N��+���nG��~�I�;,����I<�_ ��,L�W��-Z�I�)U�����ˀ�r�=.�|��QB1�v,�~)�e{Bx~���U�nnr�pH�M�x!>u�o��q72��Ռ��) '���(sA<F�#���Wв"����C���v̳V�/��x���L#�'�2���� ���u=��{-X�/|����j��X��=]��m�z�P�A�$Yzzb���`��0i�R���	��n�,���H���^Ed�~�����g'�]�w3�"�{���K�%�Ɖ�KL�',X���
q�,��#k�+O2�^uuq��/����F̈R{?�'�	B����Ù�&�tdR�QK"z�%��0�8I�m6l�|��4���2���{��7��hq���a% �h���ğ�.��-΁{���X�%�b>g�o2e1U�z���1��zH*?,q~eM��� b��(��H"��-��?;=%Cۀ��e�s{�6�jPJ�A�;��%<�-ՏE ��OҞ�-��]]~�J��F�����N�((Qu�����{�M^yI�������'v���Cm���1����KfCw
3��v����7L}��������$�\}E�5�i�v�;�=�� {��N��)���"A�ˇ�z�q��vp`���}�k��P��~��(�~���\����Ar��ʴ�t����lW�aK:���^��;m�&� BO��������!z@">�m����v�@UdúnC"�T�H���	_�1�}!��f����O�(O�n�݊u� ����#����z�u�����B��\K+��������a��;��*�!ES��}x�j3�f-���,0�$d�tK���C�r��jvj}��L:��)�(&*�5.������a#�Z�ȟ��b��dݍ�(�Ps\���h�)��&�����|W�M+����[�6X������b�H�oUu�X(����͌gݚLF�W��H[����ƿ�1Y¥�[�I�A������4q4����=�
��c�+��q(��� M0�1X��������^H�_8���J�����J��̥OQ#��d�n|Q��y��������"����颻���|)C�f�s|�҄�#�~����uv��u�����D{���#����͇���f݂��{���2� -��+���e�U�#�п���Q���7�x�[��>��z��i>����{�%br,l����ؑ���-��L�3
l�u�͡P�AHs$��b�����+��˸h�q�������T����9\*ѵpN�7`��:W��o&��q�nMd��K%��'8����^��Dv��(�(�FTTSi�P�%��%��}�'ya5�6_���G� ���tjݭk���P}S�uFG��͸��Q�� {����Ң�����ƕ�K�����d���'<�-����K:���^Hb�_	D�5�E<΄�l�)
��Y������7����ނ�{Y1WaV+
��PV��7`��t�\���~�������=�I��s0���K׭C�=�3�]q���'��G�⩦b��)� �a�j���.ߔ��I��Ȓnć�G�f60PFg��dU����S~ջ��������KtV�wT1�H��O
)6+��~�r��� �����4���J�h�â�w>\M��/���,�F��͚�f5z{����#U����°M����W+[�f0
C3���w	`�%�e�9=�{��|��G�F �u�7���G�������i��Izʏ��<2��2��]>]��+�<T*�7�op��,$���Ug>��y�+XB+����+yu��[L���ϧcc#8gj�,{%U��O��i��V������^~a1�ik�^~���!�8	��m�I�%�1���M���	��A����D�V����7�~�ݏ��{b\\���Ar�nNa��g�񅯋%5�SMѦ���*���I�s��1R��)`�w��$Y2M+���$W�he�x��F�j����Så(�2:zr��d��� I�E��]�noM~�7��l�ؕ��>8�JwÆ�q�:C| 
��E^+Da(,%Q�ǺG4�L2p)�`�j�ҺdS)��E�$���Z���@�h�r��z"��0[�D�H)X�Qν�~��𝣤PJzwN���z������D'T��}��%��2i��_�I.ɛD0U�Ĳ��M:^g.r���[eRq�;rګ�~�����O����;��nN�N��l��VY��7�%�-�<@AMߵr�2���m�一vC��Hn�c�:���s�%i�4��F�M���3Xf5F`(uë�L8�3�;E;A�T�1w�#p�q�ޣ��e�4��`T����R����s�?��JPh�aù�/�����b�l���������V��v�Ȉ�GZ�Fsה��B&��h�5���Z��&��;��ub�y�����S��T/���� +$�1�EGp�?mWp�fps���imu� ERZ���^�� �6i�G�;�I�ke�+���z�-Y��M�D|G�0��v��No%O�:��}��p����d �?\0k��{2�����e[�=���T����c�]۶IV�+5,�`�P{���OI-#H�r�a"O�	QXqn�]j�mmX:�C�-�/Le�nAv�sy?�z��M�l��$E;�G!��vn��H�{Z3c.����O�|��,&�i}�}i�ڿ��;��2gZ�Ek�Wx7gpg�	p�ψ��I{韹o�<μ3��ᨗ�P�=���NB�gY�-�� =3	`��V���'��V]�f5\{�am(C)@��ǘ@
����f���[�	�tUp������*dD��u�~ޯ�q;N=��MpM��.:0 a��ʿ����&��y)D[8�����Gܗǲ̏�%��")S\y��T+��������: ��EO�kuS���V���rص����WXʢ|�_Z�A)=L�\�xc�B{��h\�Ϻ���8���q��<5�����w��҅"�#��3����k}����.�\2l�VH�F�7OЋ7���)�΀��3b��u��}��Qz�]��T�%��!2m[i�Y�l���]�ϋ��u��U4��7d��]��Fc��o 	���}@�D��3�%o���/�"p��E���s����@�Z�*�����β��5`��q���9���ė�,���'����>ѡm��lֳ�O(�[�A0K�Kg�Mc���b�l�e������'Am�������WŬm,���g��(��,�cdڰ��ҧx�^�2���B��Y��}�y�oDȏ荾�M��c�ʭS�p�8oN3��x3����3�q7��i���K5F�l��;���J_Y��K�"e������$��]@ɿuc����	b}j	�K;�Z����%�J�#���+x٪i�O�!~��KHoG����
�+��因vn^5����#rH��^V��3clT:�`�ٵ`���]�{��$l�%�FB�����c�Rd5���N,;/�ɷc��m�W�JȚ+oqg�J����0�;T���~zȀ���q�"-W}#L�#�9�	�}ߏ'��1]����X�߿�5ݥ���/ ��%��zX�����#sh��`�Q)#"`J1�6tҥ�ooo�:*�)��f�5%s�W�k��H��SB��ū�_VHd���{@:��e�.R�,��Jt@��<�}D1�������	w���pe� 6�ڐ�����%@�e��p"�*0 �ۡf �C��&�S~��~9td~���d�xB�a�]�o
��[�xGt<��6��9����+B@ �?�@N��|�=8���'$a2����wlG���}�Q�g����q�_���IQ8�믈i�����}��׵v���	r��n�w�f�p��3���G���G&Qb rGU3e��v^ŬU#�ZԾ����vBZ̄P�#�܇��Ҭ�˘K�c2¥�ő*�(������׮��H�i��-�tRz*S"��Qji�P���n�����t�8SJ2�q���:�Z*
�g�+}K�l��|��m^�[�i�[y��R�b�= x5�����V�s�>�z��5�cGqq�g` 'CZf�_��Z�5�@�T7�fӵI��RjLq��k�k��\My����H�uIs+�:n�����(s�F�X�_gA�䕱J�CL�r�x���Z5�u���^�A� ���D��dY�lY�����'�Q�}"jmNp�B�5����]wi�Hy#A�&;ү��To-��Q���y�xÕ�mlE;���`K�\�.��%�t
@�O�Z&�]C��S�hM�@���T8i���O�×�V.V���n�_biK��L�b���6v�!����m�|����b�+��,��Z4�_��|�������:�u��(��'���MFZ=a�j��+9r{.�B��R��Չg�D�6$��yE2!��b��<���w�/8C�u?��E(9��ry�ʤ�)i�T��>�Q;�i
#�Õ��A� �K�w��k�(����!��Ҽ�k�)��ћ��UOg�<!u�Qs�X�[2%�Uţ�%׳��<eޅ+������G�,�����_�u~?��ʝH��l�����d0�qYu�r�Eh��Ș��AO׭f^�ץ����E��DQ�Oom�ve�7��w�����g�+�^���mU�b��BK��g>%���J�V:�{0��V[��R����|�A�J����� P� ="d��jF�׍�j�(�'���R�� ���5�͛5#µ���m�/K�7;���!�5�Ph����T�޺7�=s(��ܠ2 �̊���C�����\ø�<�����"��ab���\U�U��>�?�{R�*y'��H�������YH	]�/�����wM@�SF3;�I(�()��%mY:�D��~�\���e�λ�c��W�� �u��S=J�rDY����{_��hr�_�MS|��,��0[�8�m����>Jj��$�6��OuV��(@ݤ����V��)q�?�W��a��@.��Xe`L&��[#�bf���E�����e���@��ψ�k<&��$��;�BQ�gZ8V����5�r��u[ߑ@�\~��	��yy@��EsG�cEQ3�����Y�	����?C�{%f��V>�}G�8͐}J��n�2d+<�9�6"=�N�/�P)%ђ��d;�$����Ғ�@����: �0�霈�����r���H��|k�5��&�}j(3�x�Yה!8����x�%���'
��u3��!�$UVV&�U��;��Zx�/��#1�����1��xeo�"۹�~Š�KL�E�P
:�8@��zo��⑥7Q�0F�'�Lp�KRa���!ጙ�=�'�i�%����$/����{L���S8��gn�r��,�z�8���{)HƖh�E�䯇�6{闄�s���%�dTPĜ���W�
���H�/>�@y�#�_6�[~B�J�Hsc:ށD�y���"����Q0И8�"C��;@�tˌiX�@훯ǫш.�z�y�c�Ӥ#��Jn�rFNT�:�dG��H�H���ުALz��N<�TG��	Jh�lV=IRbgwI������O��r��RO+w~!>������Y8�l�ݹPo(`&Bmޛ�����Bd�ad&�'�~T�k������I���A��[���&�rM<OqAw��!���%����A����|�c�����}�ۚ�����tz�4D[�lyJ�v�+E�d)҆)Q?��@�P���\J�ZL�ȴ�0Qiz���Ǵ ?
��.�7��Q��ԗ��iΪ�o��/$�t�8���$����8�C��f]l8���{@Ԇi��� ����Qx��橌[�ԣ�뎑&E�tV���@��g��&{2E�\?�T���j���d<� �oO}S\�O�}����]����B�����Ϊ�&aQ�B����Ñ���ҙgl�|$*�iT�W	#�clL���)ʨ'<<G0����=u�S}���(�A�Tל���D���a�WU�[�K�>zջ�H�Bӎ�+S(��cg��`�q�CB����c�O�׵�@ݍ��A6Q�`� ��k��V;�9��u�o��h����'�T�8�p��t�أT������p��*�UŘ�,6�
z1�H�tV�V���<��_jBVT")���F�x���?�X�*a�>���w�U-���m����'j��Q�A�c±SYȉJ�(�=Lߧ�2���YA�JY�g�#���ӻ!4�d�&�������O7�����
j:Dn�ꪦi�m�w�_!�yI5u�@�1��]�(��Up"Q(�qp�ƻ�XժU7\d�J���S�W��a`cyḅt�+�&9#�t��|�nWE�`���ϐ�md��o������w�;ɇ>}SGx�q��-�?9���6��N�q�_)�����,(� �DA�C�ћ�Lr��Yf痆m�8!»���9�E"��є���i*Gi7��r4`�:��J�c�qV�GV�7�l��;}��������`�oݳ�bg`��{�D��S�����GVc�V#E�����Z�������ŵc�`��YS�r��ywG����a�>J̌��p6S�4���}BrF��y�Y�?�l��� &!���cjS2�.��b�]:Ղݟ-T5����-uo�Qv�*�E>�������X-���C����W����0�����8d��S��{ e�#6LUl��j�t,�7ʽ�rYo�<�u����+��*�� ��d�8����n��7(
�!.ԓ�S�_0�E/C�h�&�����v��4�[�NC;��+� �/aF/g-��턎���T���2�A����eԁ�t���{�|V���k�4	wl4����B]�y��/����Uz)g7H��yQ* ���C����p��ہ����K�V�V�����}������w�/��2��}"�	3����C��'�B��I�=��%��<)�r�JtW�{�ح$3ݯ��p�+����R�����-�F�s�����賨�[F;�;�Ō k^��&�\pM8�z{k8��b�CA��A�a�C0�4'q����E��%�vͫ�g*�_�5b�;0w�^�ʄd{�J�:+0�b�4�r�}5z��H�:ӨɨΜqu��O/�V�l���'[����TZBj/":ck���2WTLUWЮ-�~�q�j�%��oۚ1}}L��u��Ϗ�����G�&���p�R��-�7&�-���� GW�*7�C�
�ڡL&��ҖF�h��/W���v0�T���o=ޠ�#1��_x��+5�]�+o܃ja��;�v�6f�_�\9=R�a&�� 1c+ms�h����G�<����I���@6�Z�p��c�4�Kc�\!�����Ķ]�M5�4�S�C�[ƹ2��ӄ������*1�����}�ݧ�\9��#s=�����g==8vJ�]���B�j8bE��΁f_�eH=�f�\m2���t�yy��2AD�]z�n��sV9���b�� n�,�c�{o�V��%IRs��q�z^h]֋n\ӗ��kӿGNS��.O�r٢fL����,]���U���M3���ޗ�аJ�9g�ڟ��^,2��m ��6H�]Y̥`�F��v�]zrq/zƵ���M~/��QӏFγBN��Mk�y#���q���J��>�4ko�*��։ό����I6���b�`W;r��7�l@R"�� աH\�{����#�1A�Н̧�ON�ʓ�/�R���7��@�t�����7h�'hfye骉 ���4����j��� �-Įz��`Ҹ�˟U!M�d%Ֆզ� tMsOr<)�sY`���5�������e��� �f^���=>V!�,�K&o+���L[��̓�	��&��B)������_�(1�r�$�ڇ�;8ZLox���x��5�V��M�a��ܶ��`�g��Ú��>w�v�E, o��$S��
��(���O�̾��]/b���K
������g���:��$B����J�W\f^����8�J�T��9�_�N���B���-�9���W��>zh��?�҄Y����am�z���ژ,�^��C{�!WP��~��N����f�Y�Q�v:�k �� ��`Y!���?������i��H-"�ե�ސ��t�ǎ\��bĀh�Mɹ-Y�s�����DgL�����̿�3�؎{�8�B�%Ԝ$n�(�ٸ+��X��@J6&�H��
�g�ITCa���2��3Vf&qyۆ��D�
���6��2z�['��qGWY�e�`�x�i>=�^MF�V��#��:�eM��5�̐��9��'`w�yΔ�����K�]�L��_��D���?9^��q��pn� ��͂	 ���A(�$�d.b��);e�c�ǜ�*����?�R��N`�l+��BB���W���\�T%�s�j�{#��l������6�9��( t����E:��rS������i�"Ac��c�T�8V�B����۩���\����(�ǟ !�@C�n(��0�rk�Ro����GC�'��34I�d�7z7oM��ă�k�șzcM�ُ����=r�WM��dr��Dɝ:�>HK�kE�И��aU�����]g�c�0��]����5(-gr07��-�����Q��QӲ�9"D�m��}k)�O�CRs�JV֒3�F��䊔�Cl���\�X��A�1ޔ�ї8�Ό��m1֯p�����\X�Z�)f�5hl�+Q��оd�&{#�h%^�mI�W�(�D}vq�l_l����c�_��2�� ��: V�nsRbM��J[u��#��	�eZJF���D,�{�U
Z\	J��l{.���kH�0qdM������[��vB{4��$�����!p��*V�ܑ!���]��7ڤw��K��M��(�S�Oi��B؋ׇ��6��E�������)pQZCR�d���4 �h���}ςB�浸�-��I:�x�y!�ε|�|����x�Q��6�i�uS 1����Tg24�G6"x�ۇb��5
�i�c0�ɤ����:�L3�Sen.Ӂ>N�	(w�hs�����k�C��4i�^)~|l���8�m����^�,�RY��w&�;*������J&��HX:�rc|��y���n�*��c҇�R�=����
׸x��/D�>Ή��ۢ�fp[ɓ�o�!�����J�!-?�b� �YQ��V���[�F��[b�V]��*���{��9�m���͵�c�D�kV�d�U��L������}�ݟդ>����Ґ���_E�	�G�*�������~��WOF�K,�����H���ҥ���Xӛ��!�����9��T�5�*������qRp�(O]�0K����w��P������f���s�Z��}W����ۮ��R���K�N)���mR�n�˞SDi���� ��"��F9iVN�s�rF�}��Ū���xR�aF����z�p��قo�����b%لC����2�� ���X�� ��ZN��z����6X/|�|`)��{X�ʖ @:$|��@d4�b��g����]V�Bђ�^:@�,0��/��땍�G���J牲�DC\i/�����t�qB��f��c%�c{���x�\b?,�"f���:��&�S�Y���~Dٯ�Y���O����>��"a�a��e�=����Rw�����a6uFP!Nh���g#3��4�.oAB��UwƖI�ZK�����G�*5S	dL��u* 5� c1�,],�_L_e	8-��N��ԣ��P�,���Ӻ�>�c�16�cJ�i�hG0� 0�!�?�g48�t��[��o�p�[���B�-�Lv��p�O Ի�S�>ӛS<NPe�9_�MFC��^���\��>�[O��!]z\$r�Dw��x�z�F<�>��Pj~;o�������u��]����3�f��� 9BYt?X� fS���g����Msc줰4່4¢�f�0�]l������FrA�kB��f�P bc��tj1oۯ
��Z���St��1�l�3Y�>��Ed�,�����!�%�^�[��,x�o�kV��r^�D�����Ik8Y(o1W|Nƙeٺ��,�v�2���1ZŵL�1����qY�bF�*T˖�E���j߱V�'u�"����hk��m�'���:�"4�>w��hۥl�5�`aB����źM�J�/Ć���a9��w�}���n��`���2��4�յa�yR�����ߗb��оxR�Ԥ��F���������5X�*C�$)��#LS�܆^�h_�M��9N���n�t�Q�*<��.f�Oq���c{��j����Y_$��Tz~��7a��3MR�W*�ֈ�:}:5�P����R��\�u��rG�Q�����U���ɨ�w�T��0d�����4����$|X��y�|J�3ek�'��wC�7Nj�pd�ˊ�<@AISI0����:`��}f3��;7����Fݨ�G�U��V��Q��2��~dq�w���������r���Gw�g��^��ۗYVn�'̮�S���J��s��C��yͫ
�V�g�c�IP�K���pUd������˻١�>���
\�X��>��[7�u&��7c��_�8c�?L-J���(�=� �r���k����J.v���{�	��L|v�A=k�@�耔�T6ؾH/0t/=}W�]�N���㛆��{�!�i�0ua#��.C�I��N��u	m�E���X� �G[�-��������t�nJ(7����������+[O��.+[-P����� ��S�D���Jg���>q�g�����4ڜ��EhK(��x��;Ǟ\r���谝�z0Y���,��..���� z���Mocs9S�Zl���Ƀ��v�|��܂>���96hK�=PL�.�Y�r0_��*��1̲ۙL��T������Y��� ����@8,�N��f��̰���IM�L8{�2�m������x�)Y��e�Gv���1�VOW?�͜l:�(>E�R�X�q9L=P�����<-6o������u�E���qM�ե�&HP�dWK��s%Sz� �!y3M{{��oR�Q+�T�X���z�t�M�U[j~
�ҽ���k�,W�]%���v�"^qќg�[G��K�O�c�/D�N�}}v7�h��G��L�ٵA� ���q�!V��4l�y�OM�|�q�5a۠�qVǝ/���H�w�-YϞ5`��_L�z��F���M'���+��{�"zS�"��[�rD���������3��R �e��}��0wGjHׯ�oOڴa�Ѐ��S�o��}T�7Ҧ�Z�m�E@p}C���q�v�h�R���Ŋez��T ���^G�xtExzo�d�G�v��'��j�en�]FՀ�o����Zf[�|5P�C'r[��`�0)�o�۹L�6M^��!�����}B�	�Z���?�Qs��!������c1*Q�-�~����.�fl2��S.�<��*�B�w+@PNғ���Bp�gr�� �]�u��}2i���k�Xĉ��T�@�G,1S��e'z:��Ԁ��E���g��=��#�-�1�Z��:���-ϫ�}�������:��ը|�_�ń��AS�M�Der��%�+6�an���sW9��j���E�b��B��*ҌR����X���
��>\�:�B̜���]�t�TB��M�Y������<�������pDhsMgz�83���i,q뽛��
xXm���N�#ɔ�����e[2�D"[ix�!*�ǜYCx�w�[�LY��U��Y�&'D	.�u��S��-ڵ�2��$%�_n2��'f:,����J\��5�R���g���0F$��h���=@���UϠV����m�]��+��l����lw��	1��m�+�2�YG��U���9-"B��p�`A�mJ��1m�����o�v�V��X��($�lQC�m?�j%_�S��?!�b!b�;�CJ0k��Ka8�|�^��ZD��63]�;�i@S5LF!y�|Ȱ�4`��N_��/�@��oi����'� G[����2������D��l����i�0r���A��xUm�8�����pA�_�b�m�,�rQ�F���֯a���L��(��+��
Y62��T�!�<�F�D����G�Y~���=�p�n���HyE].���Ѧ�l*t�#个^\��D�*3	���,;.K�W��+8�8��oy0ބ���ً\��C=+F7����NNa;�%ö����Tw2ڈ�i�ަ����#=��fy
4i��$���a��;ǚ�<�g��^+�[]��B,��+ ���f0n!�E{2���*�&U�I� ��)��[{)�����h����J�:�3	kb���6�#�%��Y���r\O�W!��k.en'N ����ʯ=Q]�j�A�\���B�Cn�ʑ��\i������3��1i���2��$�]��ݍ�����s�W9���<��E�j�Yz��)>�&�`���mz�t��9�@��@�����ө�C,���Ey۾FvY�흇��z�E��A�m�jI��7���過����*oR��Z��d��u�=���V�� Y���7ɖ25��Y��va��DS�R[���i�T���iO��a�7W�ϔ���?���05����7��̍�`�/ў"��0�'�w.L��l��� �_�j@Zp�p��^�AF!�B�<�UH�L��Fh��;W�LՏ�2�Xh�u��B�x�I��l�n�d 0�śO�T�CC?T�Mfn>'"�
ܯ
����g�	�ƺ1�uY�o����+2�< L*`'�Ӫ?W���f����D^-��}��*w�*���v��m��ҫ�%@�DvĜy��`9e�J&�����p=o�4:�"�:xۋ6�I��I�������������9�,���(�8�m��
1�������y=&����R��V�W����W� 堺P2����=a���#������ٴ��#g�o��L�N0�[����S��1�P�|,E4K(E3�k����n�1w�E+ {�f(U��uq�r���z@(���~��V/~���6��M���޺�%?0��Įʞ�����cݮ��t�6��FU��zz��mz�q��Ƅ�����!�Ɲ.<(r;jn���`�e���[��E�S�g�����}�n=�\���g��8����+s!��-#�og�=�#���l��cΤ<�w׀���2�*���A�Q1ӵW�A�!
=�G#��W5�����`/<_f'a����$~���W��6hlt���G�2#�%K��Ș��t}��.*�\ε�[���g�b-+��]�Fõ]nT��f`���y�&���ϵ�^��z�2���6��V�O�FU�f2??�"kf݀�K��.X`�SL�_C�O&�Q)K��BO��k�\+Mث��uMT�zh_i��@M�d�!b�#ת����QtX��sD9;ї.���H��5B�)n�eˬ�w3w�]�T��J]d�	��6!��d�ZK-�5��b�f��吸	��s��aE�y6�1���K�ȇ���k>�*
�̺)Hg�Z�1�pS/��}4����9@���n�ĵg��;sK�����2�x���ev���)P{XM[[���*:n�z�XT+��+\�\q��Rc�eG0����^@G�"~����N������rg:Z"� �8��pفnsJ�+;�.:`�YV��D�__�T��hʯ4����g��J+%�F�4���z��;�(��p�/ S⩉F���ҫ��%����Ґ����b#� ㄄G�&X�r}Ⱦ;[�8���%������,h�2�mNheu�/N
���~�.�D@�`�����3.0;`*��G��-�.y{m!w�<`" 0.d�G��t��wi$,�92Q��Z��1պl�{lƸ�@�[+�%	ωW���&��m�;l;�#��0�3��OC�����?���Jw/�re��}����[�E�����l5]�+ ��9h�/�m�p_L@8���H�߆�\3�I,��6��;��z�a���U���9��̺�Pl4V��v��{Y�"/�C[��<�%_E&�����b�P��1��hoeH�~����K~N/؂"����tC�K�'�%�)����P�Y�f�G�z�>o衻�
E0a��a��DE� @�>��~��#`�Ӂ9=��e�?k0���~�Q�����]9���M�V�hI���?"->��)�� &��.���#oS��%���)pY�.}I��++߼���7̵؞��Q�%��r����C���"��١_�"MV�*$�?�i
���z������Ó\���),v��<S���JQu����V��.�DZ���/�8��~#\|_�퉥�&�\�E�� �B�A�m���*�>�:��V	�%�_T���{�Y}x=u�3�)���S��U��@����A�
�:�hk���D캭�:�ʜ�S�xP��ܵ��:]��,�M�eJ3]Yp;7]�<�r̶k �,ڎ���^�ӈ\_;eu.>��h���b��}���rJ����Ls� s���M&�T��$%��ݶ�m�TH0�L�"��÷1)^2����s���pW���I�$�Կ�P[�>�lT����L��aQ�r��ˍԂ��r���i�.��jo�L]�P��bf��;WUަ5,9�h"�/��j�kocnT����̗����qw���Us�|6�(l����h����|X�Kq�
!ξ~d�#�b�CxR���C���ߪ��ldQʯA���Gʴ��ql-@�Y��,���y��X�^7�`P.�%vQ^�ahB���(�\����ȁ(����+ZZ~��g܂.՜�f����r�m�Z��Cݛn �x����=�~:"&��k����	s0��_1�ȏV��=ٻ#E��� �{'�mD:#}N�R ���B䆙w�\��Ll��o��1��MW���B�'��EF�&� &��[=GK7°�����ie¼0:��r�&�7suP I� �����g���e�q
��G���p��%K��ͯ2��0�4w��m��w�^5�ѽ����y�7~Jm5� �Z`�{�-b�׏���+c�A����)�NY�y��⩬9hJ��}�\��È�:�8_�ҥA�t"%���K���/��]��r��T	{S��(
�l5�q�}cPW��!Y$\<6�^���g$G�4�#-��?~���3����P��6��w]xFYa�K}~�������q§-�h�{i���5W0?R���ulr��8��F��4�9��)٣@�OՇ��4����E��.fnH�RU���w�'>��>D�����w�h�,ס�_n7�o��X�f������8��F�r�Cϵ��/5*��q�{O�뼕x�*�%��qm����S��B�j�3�cjcz���Xp*b|B�jY�=�R��mհ�ڣ�Z��Jn����9�J6#�T� !:t_��p�,{A%3`|D�\��IZ��������>��ɐ��?m+�m�@,��č��*������ r_������u �u����Aeh1����U֥cz��19�8��E��e���v���9	=>ի�xeu=FF�=�0J�Sf�]V�����Yr���geI_���N�'��4�*���2�@�z4���QD��aΞ�J+������hIF��'4Q��c��j[|!h8�����3g
��{*_��;�a���£u��d�h�7���	!I���1�סu�f��/M�1���0 z5�����]� xf9q�����s�S��7�~T������h�`��Q�G{x_�f�UcS�:<��}��Xޅ��k��ʻ.1�1�������#�X��p�|�emL���y^�4݃�}S0CZp�L��si@\@��J=�5
����������!}��j��T{ǟҒ*��l�&�V论Q6��;lV��,���zo H��iW��4��t�	��Rƅd9�$k*�c�[ ��ǭ�$����Φ��g͂�A5fd�������v5 M��<���r1��r�q�5�U��жO�r�_d�s�V�ǿ��=�Ҹ����N��E4<3sۜ?�͞+Ͳ�rs��oN}8M��H�*��dT�[���XD^�w�y@8+%R]���Ԏ�Z���x�F<��DB��$�m�*�2|'pa�"@�1�� ����܋�*%��~����K,{L�8#L|��N�P�������6��ş����M6���n��`�ή�Zoz�������^��{YU��o��o%�c N���%SF,ւ���V,6T�y�Ĺ|�yϯ�� !(��?p-SCGO>|��ͦ�	Q����Z��7�h�<^�tDft�dSN+ѯ�9v�s���FOn�+l>��ag.�}��3�{?KW!d���L��ʪ4ۑ�	�;�(j{���� e*�UY��H@�;�Gr���\˴iͨNn����$p�<kL���C@I�l|�V|Wh��X5�5��o�%g���Tr��tr��	Q�\< �Qip�g�~o���\�[M��N���+���/>�
��4�hj�!>�׷B/��3�����}�\�����DVdr�p��[�dI#`��;��}���<$
nO��.U���d�(�m�~y��Csٗy\��ZR��l�I�e���O촜h�QvN�e��V{\4`(F����a[�j��a�Fb(p,��r<3�I����o��ᘒ��Y�"�L�L�]8�7�V	�a@°e+����]c��7Z)|��o���ە�EM&������*�2�C�gk�"��vtI8��,bSJg�jr�p��p~���K&��aTbZ�� �ӕ�2�}�y�ں�������6���������(B���
L��H(颪51=ܿ�k�^��{���ٯ�~��j��a��UӅ��.�PE@�D`&���Mf8�j0?�2$ �bP�o��2����c2/�J+E�w����5a?e�H���_�u��k��l�����q@��/�E�sɨ��Z=A�0��(�^NG�+h��L�^�W5���ˀr��[v��r�6d�8 H��Йt��@�{n���S�޺�a(I�\
�Q|��М���?�~DP쯡�nJ��A!{?����^-�wWH��Ty��"L�(���I�_\����mp�t��@3"mtWuB�!7ׇ�GU򌃃�0z�,4��?��@}�, �3�|k��c�з���_�I���4�Ю�mlP}���JnZp��y����tF!S���LP����?�C���7� ����C!�� ,G_j쇠~u\m�p�Ԥ*���n\(o�i�e����H��� ށ�,���;�i��B!�pʹ���	��aބh��A��`I�e�I-jq��ߋ!P�(�4O|��6}6�j�h���+�-��!A���J9ړ��c��zg&[�O�B� ld%�@r�룝i�<�JI��ؖ`Q7r��Z�����N��1;�բ�>�w��*��%�C)0r�F��
�Ǡ���N�{x�J�N�?��vM�]Ћ�C����~;)u�������ޏS�?��Y<�#�&�G�bd�mR�M��k��9S���M�V1��j,�9�V>��l�3��**�N�i�]3~�+*�}���8�e���R�tiԲ�i rWG��b���Mw�%`��|y�p�LV�x����T�L��1�9��ר���a���)����lkb��P�d���m��}c�P���H���L԰�d�W �hT��f���� X�"���� �&�L�;W���#� r���,a��|C��}�k��)x=�<Ų���伾�$�R����y�i�j��YTqc���5�N�c�{�e��i�	�J'6��������X� ��7�����B7���[�(K��[V���,���q4�B�_��gZ_�`�~?xU~��M*1�>�+/� �.�'�Pv��`�]^nw]�u|[m�g@��x2I��_ZJ��sJ�2H���3D�+V��@�N�Τ�`��Rl�ަ�n| ��2̇���I˳�`
��ϻ�FH4�PL�����٣�	���T%Z�Wj���nJ����E`&W��kF�q��b4:�h?�gs<r=�`�B�̗�O�ȷ5"��-��Q%�h�Fe<��X'��;�n[�
���N�"F�x���b��o�!$�*m�z�X۪ʆ-��(�r�W�Ro(�Fs��(,iׅ-��U�\?^5Kv/ʪ�p�O������ᆚJ��i��?���N��q@���ή���"*.�AX50e?��W6@�n�aD�,$�z�K�G�) ����j���HG���}'� O��V�DZ���yɌ �p�&�����-��a�-C��+"��<�T�YP�d1�ÿ����w�Ɗ��je�+ެ��B~Tx�����#����,�l V�^�AaW>mZgC75��F�E���TB�^�]Vľ��-,`W,gM'������d�!�L_�q�,��~i�2Q�"i�-��}��
h0�1�t@���J�\��Ï���j�z����/�?�w,�"��MV+��P�vqĆK�X�2w��qޮ��8ꪇ9�DH��i��;ܤ���2tX���S/�R��\�3�N����xn��S�tB�A�C�����!|�i�/�5��%D2�Lw�����,[��-F[>3Iz��T�s�5[��ױQ����@أ��D�N���,��}�~'@�H7��m2�Z�!��}ǋ3F�+��l�`i�.��T'��h8�|�����W�D�E��1�}Lp)>uV�����^���!k�ߔz��0����ol�,���<91f�f{�U�R.<_�5��-�.A��
$_�8[w}R
5zm>�1�Ok�Dg5]���B�-y �"��i�����sy��u�(b$��ǽ���!]y;# X�d74�s��[ћ=a�{���nBH��B,��]�w�K�NX��E���.��Ȉ��]�C��Y�&��݌�"������M�*v���S�}	�4CT�͋*Nҳ�m�ҪB=?�Bچ&�`j}��m1Q��k$�8��ǤRМ�o'�����=����]��!�{/Z�����Q����i�	+�On(n��������-��`q�>�b�!�y�*-qᩐD���%���s�ۇ��ղ�;�d=yO��i����ac�E!�{7�����Y,�'���S�}{S�F�$]����D�nb�^X�5CT���lXx-vx���I��0�R=P\��v�ʊ�HG��S7ND��;R,��cH�e�q�S�i/'\	���[�8-�w��n�e�g�C�&�����f��7WJ�w08��!�4:A T�˵2������n�|yE%aRj��Ó�k6��+Q7�����r�]-���ϸ��}0|�#�2�Q1�|&Z�Z2$�Q������W�h�T�`'�7�ӗ×Fڐ��ՋM5{���u�ѿ)��&U�Ґ_N��du��?R7��L�H��tI�E����,�����>ٵ�ɧp�ɹ[�x"A)�"?<�Q�c/�ۇ3����b|7xT���/��x�g8��,H.�ȧ�t�����J��/�z��3=�Bd�T���T�0F�!�����T��פy�;��Ckp�	#~'w*�c;N/N`RZ���sׁbPj��T�L���=�#ү���>��	������r�R����T-^u���iZj�������CzA���CIRgr��k}��H��4��f�& '��2雞��R���`�&r�V�3 6Y1Q��bv;d�Ԏ����՘I�um�<�<��q	Ή�(#ĥ��ѕ��n��p��6��5Ѐ��ܣI�G�$�"����x��kv���f��e�22}�`夭?���Q�x Ded5�S���Fqň�\�1N�? 3��6D3%���ols��Y)="���bޔ��0E\�J	Tz�#7|ȁ��J��ڿ$�G�4�U��V(�Q�>5(�E�<�]�x�\�;h(�^��ЇG�z���t��{���Z���R��l��Ӈ���Aoێz��Y�tKM��4�ѿ`��|�4�L��?2�>ϱ�"7|��!	��y�2��5�Iq�rD���)8����P��9��R�i���S�.##�k���)?�R���@hc&��6����h,aTxHC�+D6� љ?P�jX�,G�_�a�j��{���nTS��.Q싖7d��x#�5���"{��GWr����'}�N1�_p�
E��]��p��8޴Rw�g�"Q�^�}A<r�"e�ck�ր��������*�-
J��m�'%4��%����{��=��ո���E��2������s������=w��gV�M������L�S��+#t���-���<�&�U��V�64(UX��1�Z���2׺���y��!A&o�N�_��?�K�N
�Q%S����`��H�`��x��r��^�(h.Uu2���":���
Pt!`�ӱS�c��$m��p��t���t�|�Vs��s�Z^�(0a.E����-wh=M��ޢ�4����}0�u�Z���Y�.�mX�j ��z?\�j��r�eo��!����f 5Ş��r|�)�Sr�SUؕyr#]��H�i|�},�.�Ån��`�Y�b�:Cx�Hd���n��l��7�IKg�ڣ�]b4��*a�����V�?�l�WS֓�R��>�@HG��O���{�����?��_�?hPT�a��7�c5�8N��',<�m�L^�u:����}Á�S�b�!:|���%����@��g���H��.��{,�>��h���`�s��`����&Ѿ�c���}I��@���g��]��,��5<w~[D�%P5D5rds[u�� �R2��U	���a�q��Ŕ�����BeZ��0ޱ��e�d2 ��5�J�I(��:�=�?5����}k�wA��m�w5F_��^hK&qt׎��$��|��ж�s��&t��{���8�[]xOy%��/M�,�	#?_�YJ���í�_n�����:MS�����vӉ��0Q}U�v����N�O]�y,���dGu��/d��1%1��g. ���O#��>�^�����p�ls߮�:\[IM璫���Z6�J�?��|H�p�=����mR"ώ��W�bx@\�^3��}jO��ke�����]H��I
"�߈1��M���\��#�'�2Ґ��;qdM��X5��}�C�9�f�	�m��L�Au;2���$�7M�뒮�vUQ&���t>i�W�U]%�}D6��ګį !�1�xwS�#�vK����g'���|9�aց�a�q`�ȣ}�llr��0�\Hk�*�&E��5��y"��LѺ֊���U�r�f ��0�H�dFn�}�9��vP;̜%Q�-=��e��I�
����
��e��	z��K�r!u��\�����?��~!6�`m���rJ)zAȳ��x}�?}�W�?49����O,栃��f��2L�*�;�>�ť|���Z-�;T<M�ԫ ت,H�Z%��a�('�g�û��Wg'�~�����M�u���r�p
FZ�����D�Y2�R�)*�JkU�>��IiDm�pn���q0t��~��-�,_�h��J����jP)�E<�_{zD�5Z?�Jq��/�Ul���0c��N�� h�݉��e%��үo�}�����ʦ��O��MM�ʡ�4�g�ً_�"�M�l��Zn�?�`�
�˟�
��,�}u[���\\pě����c��A�!��v�E���&W�jx=H3�#���Æ�XǊ
�@�=����i�d_���:�M�F�X�"��8RdخRC���|fL;�Ds��e�N���ҝi���,�"<�K��g�f�1�;t����{U�E�ҽ��G��Fߐ/��\�V�	��ƴ�\H^7àf0n�q�#��vBN2W�]��~:�Vs���'M�a�~�(�H�
��'Ny��Gɾ�W|HF����~{��F˩�y���c���{_�<B�.X�u��ڮb�*YƩ�;�����=���BI��B2A>o}��C) '��/�[!�#��C�`��~�W��dZ�
�>S}*x>�rJ��m��"@L�6g�4�l@��[w�G�{��r'w�RĊe]��`��l��C��B-�}l1�)�m%���2�/U���u���+؎�@p�˥�y�3��5�������
\4�j�3��T'旉�����3�Q���8R5����CȵΊR�`lQ�/�%$��T���hz>l!s-?ur5��jy���C�Q�k��R
q~��#� ��?��ww����W�"���j�@�������B�_��D��K��0S���_0w���U�~TJ4��>�ϣ�E)Ґ��p��� ���F�ڒ��90��}��5���n�He����cI`�^S�{>?���Y�9����v�"*v�n��+$�W��6\A�3�/#���9�pԵ{��d36�Y��M������3�X�Q���Z�J��}U��="Y4FNuF%v��}��Ӥ�e�V7�����6��WP�
{����up��o�J��~����_��hx��&�q�7��ߖ~��ѳj�U��=��(|`1�	�̵����~%~,��?l�X�������x�X���cJ���/+�(� G�E!���حI��ڎyZ�o�RiU~ób�����f��:���Bh��kXZh�?0�����Ҕ	/A�T��*�j4m���WH'8��jخ�)��{�O���4��0�����~��.�-d|��|ߪ�'gU$�'f���Lpm.���!���K���Y��A�U���?���&1�v��
��{CH'1ʇ\mM��]t��u2�b�� d��{MÜ����{<ت(�է��P�mJ�*N�Y�)4_bP��*b�����ӓ�^6���>Lq�^c8'�+����M�xSo�x��[3�������,� ��NJ}й����8��ս����Os�݁�3�۱�Fknf��w�U$��/Bs���c����P�4��~:���!�ܬ d���nn����fe\��,Ě��d�?2C��%f-_���
G�ӤǡuQGpp��-d ��������½��'���>+���uY*���N�Y�'åG\U�{���/u�*�e�W���n��` FnG��2�;�Z]��Mb�?!�N /��f�' �q\�5Һ���~�|��Ķ�I�{Fg��/�I�͝�Ͻ˂TP�Qc`�u�6���%דY�>)�>�c�ൡ�&S ASY��2���-��'d��X���kC��Yy�=��-����
���Q؃/Ғ!g5z�p�}��#5׈v�E����\�p��1��8s�������AR��m��P2�.)�;	x_Fq�Ʋm;��J�uÂ>o���REK��tV�9�Q]���9�:�v���|��j)�����x������-�(3"�Ee}xw4r��!�:�#[/�x��\��7���ǅ�{�y�7*8�v�����'_&F�7 ^� O���K��-Q�d� D C���Sq^��q�*v��v��HP	���p�f�L=jg�1��@�.f�c�w��4*x�ҩ?Ҏ�b#\Ѿ�#�VN��vp�۫~��e�[$���6J� ]��h�S].�T�<JG=2%9HA����_�?�DZ�U�5�M!>��2�*į�ݘ5���{�P/�vp��I�`�hK�hɤ��`8���e�n���Muh;�$ 5�nԹں�u��||�b����ӼǷ��',F,[ƟԞ�N�w����6!w9|f��~��8we�\���D�u�q/�t�L�%V,Z���C�Bej��]��,w��/�� �=�P���9X��ʘ��)�9�rf��������u�D��^��Gr�~��ɚ,�H�Bƙ��4vt�eվOy����D���M�!��Yv�;�@�,��8ءc���=�O�Ѭ�m�K�E4W�����j����v����W�a�R̙U�v;N@4K�l�Ϛ�~�Q�|ي�<��u��(4�FVc�k%y��Go�OoO�*dFͦ4��M�����L�� �_���ӂ!kkx�G��M���d$=�_��rT�`����]���'1�pX/��jDZk��ؘO��)�ApZ]��l�gtN�Ztz�@�?0sB�T5�Xm���1��>�B�-za8�(h:��#�:���~�h. @������Af�WZqci��D�9�»����e��
Z�|%��̂��{�s̍�������=\������iU3��gw�:�?+��(��u�[dkw�j����O��&�Y�����$����6��X�"B(��z�Ѐ��<S�.Hs����>�d��������R�,zY	���#)6c�L;m��o�LF2%L�=~34��(�\@�>�q-��p��%̒��&+��w�7Gw���`��V��%�本0}�ꀶ;��5~���[������J#�ޮ	�mD�c��?�'��������7���Ppz��������n�̞⠖��3C`yA�嗝�(�Y����d��&���|h��4�����B����� Q���q����r����)a1�hz�@�?,���fp���������u��-1�t?��{Al>���G�4���Ph���m쩑��X��!���q��)x�T�O��g�c�Egk��*7����OǂO�X���zǭC;�}_��GX�mf���@�D	�0����O<|��(�/>�z@B3��!rw�I$�]u�ܐ����4�O���{�VZx���ej\�DxA��A"!p�a0�L� ZI�: 5N��a��ب��m��͇���V��/����j�����۟���ì�A�|e|��x�S�#qo?]y��ńl�T�W788P�
���d�X�[{��8f�}̏����2���t�2~�����ҝV�����rZ w5_�~��z�A�2!&r�x\�@1Gp�C8�a9�i{zdZ��4f����rRȅ�㰙�t�oo�k�����߄��X���A�6�Ō�Ed*�~�+3���Z�3c'i��0I�Lͩ9it!��6�	P�\c쾰x����"�@|FTv�K3G�c7q4�S �Nm����Q� ��'ӛ����j}BC��ͷ�K�r���/R�dЉ�pEj ^�5E�z%ǐ���~��o���%��Q+��W�����i���2)�$G���:Al�־yy^٠@oS�I��7P���5�W�4̇p����梻�85t���|�ƛ޷�J�A ����:Dp�t9I*�Ae<n:ɪ�����u{�1�?���i��H��N_ջѢG��aE�/��XM&rY��)�t��X�^���i�����u����v�:���貯��+���3��<k�����Lf�"j!��сR���+n��*�7�CkN�Էr�zι��n�� ���\:���U���7��� )�Z $�|�x�c�^7�������A��aO��R�C:xud��?2�]j�:�˦��:j>��ιqP�Ipy��U���8��ta�\y&��<���VPm7e+~ ���O�"���1�kVr*�]ת�/��aE�q���2��HՉG��ǁ�O��洗2s�6m��>km�F��Ǹ���m�n�S�e����
h,q'�Yw�؂�˾��R�$i���e �L����T��l�7�ο�l�/ �$ݍ�
4�}vּ;ɨ^m.M���)z�'���F	}u7�ב��CZ%����[t��2ۺ�1�l���z������ұ)M�v�m���k?$�+��"�N�F��Y�(hP����px�D��kJ��y	�L��M�<���b���F���3;w��]��N{����q4<�<���A!��0hv�ɋ>g悖,�M��{Gc|�OĚ*|+M�c�U1'�;k`!IT�g'��
�K�)j�e."O����6?Y�	K�9nW�cK��¶�jm2�Jh6��G��-m~�H͗��?Fe�Z$\;0�s����/�E���D�x��}�%�\/D��lMĖX~O<�O5~�B}�%���ٯ6������^C��1UEM �h�=
�AI@���ke�][�eo�Ѵy�.� ^����/�'8�h�{o��"�O��s0�lLOt�+'�6jf�pɳT�XԶ�|��s ��n˨k�fFk�I�l���u}[x0SӍJd+���,�6�W�s5�4�E�CX�Uy�@φ���i9��� O�E�Fc��P��i�%����{`�w�CW�A���j���`�'<!jo(dU�>m��cd�� ��v1����ͼ��B�[�ڟT�^��8wy�ٖBlfv{#��ŧ8�: '��/U�ĭɓ䲺����}����u��;'10*���V�6�Z��e��U��2gyB�"*��k��U8\�$��s	�k�Cq���pV��]�?��R��#D�A��!t��t!��TТxg]����m����U�řTPŸۗ�Y)mP��zn�ҨL3���)g�~t5w(� ��̂vP���4��~���!�C8M�p��d��m3���Gt�A��7�@�������-!�[4�k���S,y�ػ�to�˩!t"�� ��Gak���V��C;�h��,-��jS� �	x�����G��:(Uݙ���))��|���8sɗ�x����q���e7J�h��0O����i[��v6~��*-�W��k��g"����NEah0���!z�Q��H:َ��z�Z%$��G���c�g6�?�h�J�1�_�����}�I��@㨛��#W����a�c�j�������B�G49߱9x2ТZϢ3�Qc�4� z[���C��;:�pq�G���g��\M:\��I��8n3Đ�P[�����@eG+%AX��l-3��k�.�oܾ��ZD`tZK���}�� v�]�s�'�A8"Ԃ��������^sW�9,/moҘ/{�ˌ�sfE�5�L=�W��/^y���J��X�;���QWv��n�:v���*���9�$�"'_�� I�=�'5�p[�q`c��n��0��T�+I���i�u�S�-�C�r�wO+�0��yF�F��,�-K���3�Ϫ�)^�4*���;��s�_A��G/�^0��>����yGDʔ)��Ev�c�͘:^˥i^VB^@���B�Rl|�\�RB���}�?k]SB ���9�ӄe���t�-,J�o�����T7 �Y�l#W�p%������d�x/p%�9�T�U�<��G8]Z�C&ECMuێ�<�:���lP�l�PHP^OP��2����X r�}�#U�m�媟]e��y��L�\�o^�%gJx�7�:bJ�F��}`�^\~'�\O��:K|���W�ߔky�Z�nϺS|�1LC19�:�J����N�_�XEO�m�?u�Qfґvm��x��-�#4Ke]���5).�'��`Q:u�÷X�2�YG��V&��(�6�8��aY?T��Ak
(�q�(7��
!���m�>�C�OT�ei����ff]'K���׃��cq�"9�QswZ�M	�wh9��3�(�n?��ep�0��uO߿Y�A�C%�Nמ�hc��%���P��T�4�+夶?"�델2��6's��f-UI�Y���.�����ws5��/t�0��+P�j�zt ����EH�s�?���C�S-B�.�='�������2��w���C�����G�t}3���h�|ǔ5�v���[�[q+T�\W$�tq��q�� ��>����݊��N'�G\I���D´��g��#��#�-��k)8.C���6��յ�̃]>>�)��_�ȳ��r�:��S�����AT�I��Mg]�W�7L��o*!i�N��UH��ڬ����#8�鞃g�~�O�!�� �����Ea�tN[ g䳰+���JtT��*�o��0�W������3��׋±?�%#o�����dR
-6_�N��]�^3bL�D�"N}�����P�Qb=�/ԟ�V"��X	�ۢ��o��>�
Zn{����1�%�~�>��6w��F���|kr�k�ˬ=z�.�LPY��ԟ�ώ� 	�oؾ�&�eŊ"v6�����[� -�T��7�l�M���O�Iep���`l����h���nC2ꢞ�9��6@�c��c�2oib�������'\«*���������6N�7���85@$Mc��'�f>%��E�9|�k�n�G����c�|an�,����`,V0�����*���߼F��K��e���'�X���J��9&� m����Ͽ�F����G<T�9z�ب��~$�rC�a5�G���{�7����??+)��d}���}m�ݚk���$jr�o����A�>�:�����M��NӊZ�uAj���@~�6K ���ѧ���#��H����M���1��T"���o����cU�a�b[sеqEǔ�BA���M#o������N�O�ԳC?�o��hP���Cx I�qgK`:�h$�Q� ��;s��+\�	�Pf�9f)5����Q�O{�jCg��$e𨆶�X�$+<�pm~`.�]ܲ`)�|Q3/�h;�N�z��!�k6[Z\�l�w�@AޠU�����mo�2Y�f���Ķ�kH����)iv1�e:�9·-���O��#�6�k�^��s�}�Qͱ�2�[�w�ob��?Dgwk��*��k�U0$��'QN9V1ˌ�G��qz�7��'��e�V#-T��4�M�=GV�(��z��~7�n�Ռ���i�8tW�#(�JS��{c8ӝ��G/�Kb{�WS�Xeւ?�/\�:O�98g[�3��������ksA�����5�$["ڎ�'ϵ���W���o�:?GB=.7 	��s��	�)�[HW�T�G�f�r{����Hܜ]�����WO$�1���H�P�5���)匷��Go����Z��Zkͺ��_-G
Jir����@8` �-��aA�̯ac*�:�:��-Է ��8�k���	1������/CRW	�^R:d?'	��ڋ��%�
�z�Z��P}�b��	M}��ͤ6�	�p�rZ����JE�$A2���.��˩]��� ���]b�����ۜ�6%ng@���/�bR�}���у��II�󞬢��������=Eq��>N�0<]�#;02��=O5JEW�x��1{����<?�	�pɧė�X���B��GKb�D��j��eQ+��_8�!�P��*a�-�r�2fE,b/Ͳ��az���EF4��[D�ѣ�Dz�&�c_�y��]�~�ԛ�Մ�|�U�%�(��8�?�(�ъ�pj�ѨBѡ݉7�p�s��y� [�M�G������[9&����{f������P���&���4�Ufm�o�ґ6��~-ԉĨ�;�5S�۫d���~�wD��I�y�j�C`TŘt��lj*�@�H��#�E L�\�ęI�J��}̭�w���ZU���~�`�nٺ @c�X�IZ|ݐ��QA�&�a�t��w(6�$e�����N��Z��w�Յ�nw�_����q��?�6�?�l��fu�	���9{�� {s�����i�*̐�̠h�'�>��3��P1�J�Tó+��X���BK�l��SJj�b���oG�/�_!pе|�S'�(: �E E%9�� �$4��|�� �I����|?D��1�  �YjZ��˯��.F��|r+s3�0�&��e{{�5�AUbG@"��V�T
Q `3%�˹V_piΧ��;PD���d����ҟ�	o?.e��݇R	��
|u[w���!�:^t6"+c)\#�X�iM��6�ێ����f�Jƴ������Z�F��������5��ocWl�H��q�����5�Q�^�4�S��\6���y�x�)�(? P��6����.a�P�X:���ummVD�v�'(X\���#>��duDc���Y2�{�O�4c\�D[����>`�ٲ^#��)��BW�Ԭ�a[�ǿ���Vٙw�����q'R���vY��̍u���O�����o�\�Z�.�y%�Ȅ'#�\Y��<�i��;��ϕ��Gʆ�|��a�V|�c�!�=y3L�y�K��p�y;ȆC��08ڕgm���~�>Y��lf+3�r���5�c��vjq8}��or�a�?���h'�qϋWȵAǈ0W�� xO����ɻ �L��"�>����ҝk��mS�C�	RyF:����Y,� ��{wSd�IԱR����c(��~���d�Y!fK��� d����;��������%i�X���Ȉ��U��V���	�:`5��^�Ԫ�e���v�{��	��Ǽ*�A��:\���X1ܫ1�����@�y��f�֎�9�b��i|a}��\g�&�bwy|&>@§L��x���-�M1�Rp�X�����������K<����F�t��Y�!��<�W>���r;��)��j���Z���!�P���̬*a�"��a&	RwzB��4<Ei[C.O/��x��/u��\�l/��>�P/Γ੩�[�	?������<M�3b�d�_��=��+L��5�񯦫*2I,��iy˜�'\������[��o�����P�Va� z���Z�,�Se�������	���̡���z����Q��s�b
1m��#;X���Z����6�n����N���r������aN����8���"�C[�7?<�I�L�E�6�98t��7�l��5)M�K;��Ke����?-��61��߽v�f�.X�,&2 �)�߅(�OB,����W���I���o|?�T�+��2����7�ƻ�L����/
�+z|���͇u[�Q�t�Z>���X%R��r�-��W��C1�f�sB�`�1Fϴ-"�peB�b�,��'5%`���G3W�<��:Vo$BO~�E'��n��#�q����e��a�Y�PW����	<��(B�����
����y��4��|ы��B��C�q�)T�a.]S��.-j�8��E�c�>�{&���}`b����[��<7Kl�Iq�b*�℥w���/����%�M�p�v��|�/9T��+�1�i�������P�e�d��-2V�SVk	k�ýyRD�2ĕg{��ބw���#y��^�Z���U�Ls�82R^Ҥ4���r#���!p�yS�1�(�����>��jdk�$.��}@�(h�}:�������\�{Z���{���g�˃��Y�?��Z�}=��?3��^ݤ)\3�7�j���Rɫ��Z���0M%�Њ��J�3e����0G'!�ﺄk����1�,F�$JS����N�o��ވI��@��^?x�m�yX��!�gۺ�[��[u�-&��٪$")s�ǖc�ZƁgoV}�2�|M�\�D.�v@`�Dh�Ik�mA���u�Rk@�壝�D��+FE���::�z|xyW:TJ�5˽��H���c��<0�������kuW����b�j�����+G9�C~�P��$'�O<�	�	���.~i�h��zܑ14�l�G}�US���Z���.�4�[�3K�@��OI���[�(�~0	�U��EjV�\�!�Q�� PXQ�$B���iٝ����)\�)�ب!��t#�y7>�H�`BR4i���h�@1���Bڧ����:`�>A��U�X�.ʨj�n�\�`����FY���8cm:�䛍���ɂ�����D(� |�Դ\M���(�u�-�<��vVt�V>oU�#"�����y��~e´����E3���i9ҫ�I~kd\=�[�[��"��ј��f_ڃ6A3�٣�k��a"B�����R�O�DCU�����酟�5҄�` ���1��T	���q���`�+� %�`�':ۓ�2߮��&7�֚�t�N�Q�+�N���	�����I?���K��qW������(r��3Q��*n�V�
���Q���I�`9�<HB1c����oѻ"�����	ŽY�q��YK�u��b&�6����V7<+���1�ǆ�1[A�:�cp�@��S\E��	�2�7�kv0����w1�x2"�73��r�"��t�[+4��������=�H�i��$U3���nȡ�	kPe'f]�.�O���"�$�,�����mQ����̑�fq)��1����o<���BЋ-�r�OqWE�N�@�Z֯�R �Hw��8JIO�-��v��e��u�g67݆�9p�������
�����Q������m�j���5C�rj���.����,�V�/y�"����<������<��n����r��7�A���"�*��c{�g9!|P>G̈w�@IW�{��uMD{;��=�o&��p�D����^s/��B���$�<�/i��F4F�dvjZ�U]6�ULN��~4�qa!x=t8@�� }�$<4õ�S��~�9q9�p�ہ�
*>����7�=%�_�
�!T��J�wdw�p/�p�]֭%��E����{�>��_����B�_�O	o��o$ܙ�6	U 0�1~}��� �T\�9֡r�����9���R�;r�w�?���%��d
:�����p�F�7���dmIg4��M�<�[��rN�~K���
݇���V�%��-z���B5y����F��	8"M��V)�����D)�d��颋e@;�?|�Ю;�RO��,	>��Em�;#���x��/9�C��h���	J@��z��˴3�`CĀ>B �A˂e�٭�O0Na'w�1+?Is��*r�c�����K�xE[K��D��V0y%�p�ڃRhA*�����`�5
j@m�W*��:oꬩm�*q�2���rX;��_�HQ`T,F���Q�!_��`�=�Ň��p�o���T������Bj,�0�������1�{��>���	���o��#�?�U��|�A�pb�MCE��ݙ�_Q����_��g�	������ob1��[��^=`���EQ�}�L��DeWGWZ���gyكD�E?��wOQ�h�S��e{H8�h���@dEm#�!"�$ر�c�����{XY+ئ[��C�(I�I���b*�N�/K|�onF;ߢ$��FV�"��0+��b��ͳ�|N"����˼E����#gG���0�J�1��Т�~��Xy[�"�O�j�~*l�T;������C��3_/���D��b!�g�Z����`�sah�ö�x��ˉ��v��>���}�����o�����f� �QNT�����Z���4.��N?�O�P���`�i/�%��@F=�P����e��SH?����tep���g1�&h�� H�L�i(������~����9Î$������ֻs*�\[���(6���֘�3����TW$�D���v�5�e�s���"��`�a�t� ��|�-;����%�b u���k]`�
U�Bg����%�7�E���:��Oi.��	+7շvM��(�T�rFj/Ie?�O��6���4���5�,.X߶_tjs���5�U���1�Bi��u=+X|ܬ���7�h�n�o殻A �ՙ��8*�`�j�3���E�����4�QT���|�xڑ1��k�ȌF�a�#E�0�4O80��=W�7�^5f�TYb��d6��1*�z�*��>P���@�m=�֊÷IC?��ya ��
I@�H�1俦v������b��#�j|����q���e	��"�A�̴�7���j��M��=�ゖ{��[�,�*�_��H25�!��ꙑ/�6�����{:���9DI�Mj
�]���^'צ�����K6q�5|p>���Fy�4��������n�1�O�%޺ׁ�ԓc|�/ )���Y����lG?�J��,u7�i|����[���ߴ�jp�h�%�˖O�^�є��/��Em*����:,��A���ز9_x�v�Aw*$�h5c��`����npDW5���M�h��v�r�����{ݸ��]�~臙���-l�qc��"o�`2���������T�B?z�B^�hU�^-���V�aM=5�{bB'S�(*�PS2<�0&QŲ�ṖO��Ғ��?�onN�ػΊ�#?����;UGAv�'�/	.a�p�7���x]B.�[����f��5�dfx"�C'�/�;���v��R�m7�x��n�H5�64�f��'���B���l�a����B(_�x#��ٻF�>H�����x��8RY�2�N�/I:��9�R�y�u۰:��L-��@V������}�!5����sK���%��̆Ǭpص�aaQ x���3�������dX�M �"��Hs�S7*��3�,30p��(�%�'�$9�ʖ熼��,��)�]NN�E�M>� W���r*���RV���~R���d^������m�pc 3I�eo�e�/�Y�=��\ Q�a%L�P'�ق?J��bΝ%3?.�<M��R|�"���Qh2[�N�7��S=B/���Yh~\�SL��2�ҬU��`�85�,7|#&�Hz�CۙO⃀�t<���ӋZ��E�X�%���)�g!c!<~�n�/�m��p�E1l���C��Ih�� )}]M)g�T$��LAbk��I��ڋ<�_��b�F��SN��AC���}�M!��S�✐���_�r��//��P��Qn��j6��`� �$�߷�F����0
:ŴdȆH��j�}J"�q�����P��ױ��.*0~���s�Ua��:�LZX���y���)�^R�����{�v'������s��n���-�FI�kw1��$:�B�aF�+6�~�u�W�iɪ��W�P�0���U��i�*�V�v���)^�DH�qW#@�[�*b
)ɉ"����' F�3�q�7�F��gMrj,~�:�b�X��ST*��P'�#ֻؾ�c�U�i浒e�o	��xl2�k���R0�I@'5̚�C�nA-A����O/���^<\j�X�tj�
	��hF�6����1��7V�҉s�|��υ�cz�)� �v�yv+wl�o�<���z<��;��6249�0�����N��[�a]�V���r�y���!���}���:�~��Ո?-��_��,'9��5���n����)�0g��:�/�*He=M-5���چ�t�T�	D�����\N�ȸ�MWŰ���eHu�E�s��mT��O�A�D�whF�V��#_�X��֢oł���Ě�`˞��s��w-"���*}�rd+�O̧���G�\�9���!��B@���� �{l������]7��h�복�>���_���
L����6
Ij����αڼ�D��OR�k!��N��O��V�0��Xfm�e�q(��;ꡇ�sph*2~�ۘ���b��c�"���Mq^�7�D��j�X9�F'��!q��E61LCxe	��]���!�f�+�cB[�sC�
!�jڷU���Y����dKN����Ӑ����Y7����m/� �he���A�yP�
-��<{)^���(�8�t�*Q*1,��\������(�0?!O��{*��������<��?�^����$	�t/���Ճ��.̞&����$(6��3�t4�G�B�r�;ր4S��LeQ?�d|/!=�v�^)'!��@�a��Z{f�����s4�_u��.Z����9
������@���]�J8��H��&��@ Cy�+�>h@��+��`&��1�f+�a~�p�8����I�#�0Gz��1K����u?�,��@��l稙\���Il"RU���n�^�)�Bb��)2�EW)��#ѿ�����υi��x0!R���'�G��??_a�:7ѻ��5��j&���Hpp�mB0SP��RO`t�K��Y"����H�NU WE#^��\��L\�LJdR>���i�#�#E������8�����oE-�Gh�Ʊ���ג �-]��s�2$�h��������I"�Lb,�b��MB���7�AB�[�8��\��.3-<��i��
 �Q;�n���\�����#�a��8�@��k�{%�l\��F���'��t$�m�G0ɝ����j��8�h��A���.�O���/��v2G �5��+��\l�w�����Ywk+������8.pGL�2��m�Q:ܜODYY���R��03��ũ+6b�VsA�0�����@�"� �M���4ҹ򴼙� � Cl	��+��44�DK�֍����Y��|�!|�v7M�i���+�(�s��N"�G�����UIؘ��mW~x�:��$�7�
��o�洆tv�`�w��
8�UM��|L�����i��X��"�G��i�i��ݫO��NR8W�s���<o�uq���x�|�he.=��� ����h#����x"{��H}_+�蓦,߂���d�1â��z}�L���h�+�G}ȏ�}_�l7��z,���@*����W@\�B���Q�?��{�H��|*�d�$�-�/	������xd0�ƪ�.B�7jb(c?u�4�S'5�G͖�W�pIQ����VZ��3�����nq�w`�h��F�y��F��s�Fi���V=�u`x��QAn��4�����t�2�� ����:tn�_{	U�T���_ג�@K\i��M�<7Ȋy�����ԋa���l�;L!��1w۵��[P��f�W��T� -��0���>�D=pG��¢�x�Q�����A+�k�{�Ҏ��ݘ���-��*���@��Go��~�C���z�t耭�۟Q�c��KʖX��	pʦ��%L��
�!��k0�D��啢���f�,!��~��`&��%�^�IZ�oU۵����Z���%ۿ���6[�,����+�|ﰐ ��>�S�T��=0����U��'��FS��B�yK���*�ؙ��/���	��8�w��͘n��}Hmu~w-�
�Ɠ�g"6��2��]�A@ɢ����/�*��G���qدx22h�4=�ٖ4�?�j�T���Ձd&�4Ʈ�������V.M)����Q;��c���{�(e�+�Oc������Z��N���tf��o$ ��gW���,-Av�UGlR��Ǣ��7_x��D��<G�Գ��m���-�I����w标�Ӊ���e�sM��5}�w@Uu�9.V��nL�i��kz4�<2#�T�:���5+�?���h.��!���j�BH�C|Aâ��s?\�bpE��F�µ;a�mw��X#�&(�G�����,��!�f�������W�]ҠQ3h$9~cz�� 9^T�X��g�&�U-D��8��p�؜N��2�z�-H�� ���Ԫ�XR�|��N�;��h�x�^Z��CU��I�loD�S�7�q�$�Z��1�@[�|,
��ƚ�ՐZV��Y�k�r�c�i!l��v�;>��|�w}�v!݋3�u��q���n��b��7��tQ:�5�̮��u����&q	vr�����U-Q�5u'�V>�N"��s7U����H�`I�84��ŧ��~}X7%���)�&�O��d�,���Zo�M��E&ِ�[r�z��ϝ5��Cw� ��VVB{$��#C�A�!�9Z	eX��Y?�4��[贶|6�W:1�ɥd4��J�E�\S�J5; �_����!9�[�`�PV;��h�S8C(�N�����^�Yq;~�%4��)Eg�.@��Q�`<�WǸCQI4h������p-���]0E��0v��kRlV��a�%|��9%D"RA]����a�Y��wƁ�[�"�|���f�9��ĵGX0<V*�Aw�
ʪ�)�i�aI������
�����\����<�F����Zg����i'�v�j����X�S��2������<@�2gi'��8�@�p��>�Lo\D#�a�Ӕ/�x��d%8�f?�ޔ�GMz	��xY�Fɽ�R�.A���c��)+�����C�O�F�ݿ���u���Z������,�"V���%�2� ���W�������X��p�z'�b(	�k�mF�+9��Ѓ�'=�~
��֤]�c34���8#�@��1�=p��P���r���>�X'6zȩ*�A������U�O��A��F�e�W{�|��A����J�UbS����	mb�cϰ0;�l'���]�x��F�n���7,��3��ހ[�-C ���M�o:w��$�L(J����`<^|D���.Z�T?������f6UP۟u[{d��"�X�ͼp������k��ߍ�Z��^��T�2�K�J9�d�?B;�;��|���˛ Zj�7�Kz$�$���� {Ź�^a�*?���L���e��R��oP&*��>a�԰Q0+���B۶��L��>b��*��k�1��p��ٲ��ao�xw��އY�$�+W_��/6��iU�K�t[��x�n
���cXu��K�h��/Q�`��BfByy��� SeH�/�uc� +F8���iM�X�ER_p�g��cqE҅���z_>�����ή&�d�!�!`���Ld#L��D:�ĨXȢ��bpU��CV52oF�Fu@��� ^tC���7�k��Y����¨�+|�R�ݲo��v.�~����U�*-��:1�������� o�?��L{8u�|�7����b���pʀk�Q�гC���JϺ���(F�9��.6y��t}̤����F�-W��,gj��l�\�?B
����zŦ��3	���x0� �����
�¦�P�3�ȣ��$�M^���ݢ=��(��&�?X*�#+ļ7�)Ǹ��ɂ�%��Y��AO ��%-�ڧoűXc�1?�ӣ�VYF��%1��{%� +��@!��{�/{g3;�2���B��'��*���� _>��Jɱ��8hOb��}(]YO���@v����U� �+���-*�Z�*����r���q�G��Ԫt��	����H�~��-������y ���L���Q)G�o9��QOB�b\�<�k�a���3�@������Fbeb��=�Cgt��t؀G��,��Nh���3������wblCE�A�U/�H��w���?����2pj�u�h\�n\zЇÆq�T��F��q¬͙x��؋鱢��r߻����u˘t܅UL�C�֯�^,�t{2�����o��@�3������~ޘ	�w��_�y�%����<��:���,W�@��^�����!B�\x��ֵTw�,i9ǖ�;nI��*������W�a�/z�Z���?h�����v��J�@r���@=fU��	�Y�(�&�����țݥ��իmI�M���j��v�\� ��)��Ɍq��o���������u��X~�C+�&�ul�力~X�l��w���X�fmo$��� ��b�7B�L�/&r�&*��p�6���Y�9�F�*B6�@y*�*+�ڣ���y�^���S�6x��H@?௷{%�V��i\_�f-�8+f��x���M��,ځv��B�DN_����T��%!�xe!B%�^!��w�A���[wCE����z�0Q��6P��h��5`����8	ς����").ƺX�]I�^��r��I��f�ɧ攇%T�DnK_���>t�&uҥ��ҋT���U=BT����"ܲ���?�ض�O��p��6�{f�+GO�%(Q�>hD�����m�9�W6O��u���81D�*R
��¨3��,Т��8i��r*7��F³�&L��[���0*ԡk�J���h� �}$�Gd:e��F�n����t��1�4�ҵ���5o'cl}V�\��yH��G�B��<^US����������U!9��%�3�cϏ7^�c҇Ӝ�ʺ�`$I��z\-忧p��"�h	���/7��kԛ����&������K�+��=������8� �n���)�~#<����^dQ�!X�4V�P������S��_���jV6�k�7(��V*���R� �EۤqEr�}�j\����.l�e��$�g�7�
z5 @�@xO4��I=?ͻV��⯦pcQВ��&��Y�w�����[�D_�G�EX�6��|�_HxgD�wa39a����S8�-����B�,=�&>⎕���� �Tx���{��7¿{-k�D����5ay��[;A��&"�� �oR���%�|S�  fl�)E��Z����v]8s(Ǔǜ\Wp)0t@/OҀс{F������!��K�h��萺���1�;�I[��%"���l�+��l1�N�;���Ͷ7�r^ ����H��r)��v��ٛ���6��u!dL��d���K����FR����5����'Ny+l>!c��]5V���hԮI�%v�%�h+[�ai%�y������q��/Ǝ�  _pmrn��@S8�@���%��UmHAD�!�N�������n�֦�w\�ħC���WD)+�T���_0�`����&	H+*'��Q/W��u��4��9m/Du]]z���9^VS����j�|@�@�=��݇���D�,�˕�F��[���7��[:���y��e��WK� ]��E��P�RU�0�H��Y9��
��kw>��Z��v��W��WM�7.Ss��:��Ї�mE���Q7UhwV��$5�c�Z'7��*FA�
��$4�.��U�r2�\�xu?{��>�q]���5���Ɗq�}r��ӊ1$��
��{�m�W����и�j�P�L���]?����S���1�;3R��]3��0���k1��Y��;ܯ���r?Ae�*>i�5��Ѥ�mF�|ۙ�NM[��Uy'���-�Q���$%�2�j�A��D��z ;v8��e������$;��_��7N$����xzO捌�����J7n�,�3S�0�~��9��a�_ݶ�ל�A��$��6b?b3���5��g���/�	��?���Rl�E>�]����pU�����5�a*_)�����|�O���-x"�ZR�ܕ�4ً�Y�^~��@���%4�]�}Q9���	v�uGO�G�Y	�c�'�rS��dM]�i�m�-g����z]���]�~�nW_�:�9T���K>&G�����溰<�=	b�3���@H���q ��3�F1�C��2L�ΝW�sB��c_������1����k9��m�g��G6-�3�ǝ:ϩ�+��;��%-��Q/��l�$�4'1�C�����zY��=�=�˲!�b_D���a�.�K3c��1LӤ�B<�A�5��z�Q.+e�(�GrN��ILë����]��%�Ƚta���^��Yw��o팒����NB�3�m�NƫL�u�u9��ٔ<����	��Cmd��ۊ���Ko�p~�*c�g���=+SYUǌ����S���(z��TB�ǖ��[��׉���r��A�K� b���6g,�`vU��uf����tč�k�y��IЛ[�v���0�7Ղ�a�qwM�B�g?q�}*UZ)���G�v�F���>�%�8�=���\8�V}޳�
���/i@Xo%L��r�^�E��SMW��0��B�%�5�U}�hDA%I��93z�ȷ�=Nυsz1��M7g�3}:�>ju/1GET����z��	icǂ;3ô4�4��h ���M��X�@�1�y����N���u��*��#��V��.~"{���Epv3ĩv(�����B�[A�Ef.UQ�|�Lz�tH��7���v�)�����B�ԢA� �5ir b>=�~�����I!)�H� ��#R�	�]��GJlz��ag��X 
��q���h��9d&Ț�q���V�Tik������%�	I�>�lC���-Jd#�x�S*���.LH}@P����K�&������tm��㵊���뺜*;ɿ�3�GW�L�1�0��,�~��q��R%�@`�(q6�m�W� �� FD� �a����>{6���I?U?�?��m�~^�B �������`��]FY��w���oe���韒���ο��*9���7�Ǯ�����_^,8��6x���>I]�9!����K���L#����mrqxr��� ��,9�P�E���y�;"y�ѓ?xk�}N9P|I!���P���5���A�+.�Ď���Z���.5{�`t��|\�77�"̻r̬DZ+����B�!H�S+���J�X��+w��4K��qcqB��gU^h֡�ldK�T�T�/��#Q�T�.���q�p�WY��q�j�𩦉�2_�1׺�z�w���/I�O�����{g��OX\h5�B)���2��b�k�^}���9;QgK%=O��,�gMN"�>�<8c�p���̏�`��`�=�2���Sʤ\��X|�
۽�6������9<S�vwD�Kx}X�9%�QX+����6���F_�OȆu��1�pǵ��2dF2��M�V���+�흕�O<���|��||�����9u���vD�|��ϯ#��S�"��ƊnYQ��K��?�8���d��됳`������m�%��C��a���Q�hZX�2�4�BgM,B��Sْ>8�*�&�UH�RJM��fu,rW;�I�;��h�0��J���z�MӭU5:���ǥ�����>z�o�N/#��������4
F�KTC�	,��h��������݋蔂��I|��:����d����ȫ��'�g�����^��Zk���v�����c��&^��	B!/L�F&����{0�%��Ҁ�״@��[B74�9�UK��"�g)�IM)[��.���a%�	��]���l�͑�����h��x������T��
~���k��0J��:�V�ö��B�����hJ�aP&:�zmR�ws쎪!��*s�t�����AQ��.����]�Ct�K�_�D�@�;�b�g�Uz���s�ui���	�H�=MH�������u78�ݫӿ�y�io ��5#��x�{v���N{r�x��@a������"c&����[�7?�t>-����2���}XS�73�����/I|��,*�w]΅���F�ܸ���&0�T�*Wi�\������:v�]�J�!��[`�o�3�0��kQ�i�?
�ged�au���S�KFK'�������L���	���$�'Y�gb�=β#��a���e�O�wD���^'Y�,��蹨
��A�1�!I���+�5�L���$��������RK
�s2�}����몵hf�@]�Y����#ެDq������H��sQR�=��G���.�LU�%wK��s�
�� ;�8A�W� �[����u5PGp����>��7�>E��xZEZ�p�	7U�9�i����eT0F5,븩b�ݿ	vlnc��>\�\l���Gb���.��u�����x���^�\Wf�j�����G�Ѓ��l��9&XA1lsˈ�Q"p��U�}T�U� (��<$��-s��[���*G���M���������]ТN��*,;��O�}���ZHߏ|�̀�}��ʍ������:�6������j�)�_<ɭT���P�$6�)|_�ox;c��		���7�AF���?���~}G?FL�=��B�i&��+m������C|e��@�B0H�uӼ�-/S�:���1I�0��r����Uft��5gX����~+ &'(�= ���ܜ�
�n����P��e��m�,L�e�6H����2h��\g�G�1��b؜e�mX����r-�������1U�<��XE�" VVYo�T[�5�$&���>|R1�*Z��~e�n?����n��]���ߏ0����#�����[Q�����E��mr�h�S
���xo���ٛJ
��$|�b&���xֈO�w/C�Ϟ��7��vF	xrD�3\H3�M��T[|��E�g˷)�P[��ej���nd �[t�?y���&0��2ޛd�(FZ�K�$�D�D<�bX��Q�뿷��ܠ����K9_�7+`������9?�@v!�� �����>�p�Hp�q#b��3�ƃ�����cd0�3YӞX� ���.��G����7!���8*�T�t��Z�a3 �R�RI���	�tt��3x���Ŭf��N���(��*!�CE�M��+p^�v�p���%��O0�4!}�IYJ�qSG١�)�e]���� �W2�ڗ�*Չ�dmgo��p�/ܷ|�#��`�e
T���b̎;�
pw&�X�J&�j���l ��o�jPL��p�H0@��]��,��FB]NT聳��ņ�T�e,�6�u�����54�ś)R���2E-o�n#|:����3-�Ia����<���/����J�|�e!ѦXy�ނ�#��hڿR�P\����\(��ە�E F��o�ZP�5�N�~T��ci~�[�9�`"oH���V��a�z=pS��3D�v����I�|ej�>�vXw�\��20y���N�� �	LW��V�Ɂ4P�{�O~�����ꍸ�"�Z�_�/�Q��O�VKoǆr+g�O�A�����ު�R��V#Ѡ�Up�)�#���p�!�|QyJ,=ɬ����>$E�tq� @�(��{�ƻ���#N�l�����Y�Y{�k���Xށ��I�a�Ks>�-��L\� �+Ѱ���z���#{���9	2C7��[)��z�3�r�q�A�hM�yf"��]�sʪcB��G=�Z�,��.�~��=]©3XA �v�� O9�&����u��[�}@\�����M*��!���N�4ﻧ��ǁ��X����/��2ۮ=��/6e�(�TV����h?�6~9�s}���cGU	�6���n�o\:UC[�G��!L�T���Y�,�s4z�����$�A2fQ�.�T@A���l�P��D��%[V������/��hc�Te72� �Mb�a�r��z�o�qo�x�U�炔\\e���퀡���*_�5oZ��1����6����Dj>֪������߬s��ϩ�]1�RJ��	�J@$��~��+�sn՞�����)���Ȫ�ͬ�C%9b�g�.a���j��������\���������@�TS���tcJ���&��ݼ������-A�f^�.�!S' ��;���5@0�o�v3Y�d'����w�WP�+�Z�F �䯽?/�&#�7��Ҝ��[�Q�5�UT}�t��wΕ���Ƭ��������9�0^@��-�z"��u��0{�8�|�sPX��A=�Y�y�?�q�Rj�G�ʔ�ǅ<�=�û�ɴ�iؤg��Rgmr3<� �ߠ�5���1�R�?!m� מ,�ۏ��'���늞��e~�0��D�%�������敜R�o� :��gw&߅�!�ҽ����N��`n�]^��m�>d���r.g�>ei2�ɞ��U�).!���V�n���Ϸ�oF��*<İ� c 6J7��N
�5!���+Z5̰:E����0�G�)�cUO\�9�Sԑd�Bt3P�ͥ��,�@'ؤ��r{gC�bPQqt�nF�����?Q���|C�-��D��Q�B��t�g	��Vwy���D����ux�T&4%�޽Dо^k���d�j�A)��9k��MV� j&)x`q����n�܅^��w1����c8��'?~㾢�k������W���տL @�XJ����k�;�=��A%Ur"qcC�NX� �U�N~$.����'Dۦ� OI�!��w����\�Z=�b�,��x����2����+j�S�/��>��~D=6e9 �.��x#�	Q�({�4H�&T�"��ۚ	 ��ɿ�N�x1p3�E�!&�F[��֕�V��w�{#��5[6H+���.t���U��_v&�����h��0CR:TD�_Ik(�N"���g�]7UR�H�Ic_��T�l��xu�Y��-���n�M�Hr�����q湵2j��w�
২ٯ�@��L��B��|�j��~���o����Y��¨p�g�� ���� ��M�
S(�ؽ[���eԸ��!ϝ�n��k�J�=�e�m>ǻO�<ȏ�ԙ�
�,c@ߥ�R���1��N�KX?8��>�P�"2�L�r�v�c0~��ض�F��.BN����Of�7;�[c*���
���f'�*b�צ,Ɵ�{k�� "ȵ+�g_@B��ț�����1����Q�6g�ϗ˚V�C��Fx*
�Z���ٓ4J�ܢ� 6 ����K�9��I�3��mx��i�?�V����>�=����)��r8��;AL������;���vQ
��%ÛЄ��$-0�5�A�ð���RA�X.x�����t�	��E�jL�MǤ�)�˖�R��H��曦�]��}G���F��F���l��wtan��䯆��[g ��\i��a��
�}�\��w���= �4������9m�D*���dU*��?f'u�~�l$мG��
�Xt�!6,tJ����q��$.6��#���R?�G�޵���� �z��㣟��u�a& ���+���^����"��ˌ֙�
�5x�kmP��i�5���n���$DNӪ�Z	�!�ǣ����p�6��2c���6�r��0����#UG�������ц�"��/�c�9(�[K��_�u�^��0y/��>�zP������ΧZ����n�BУk��}aQ��mF�q@���M����U)�e�@u� �1��3}#�\��d�����Qƀ�I��̳������%�v5�R���������7'\=�,v��ZG��4�x��5��������}-�HV[O��|<�LD��C������;�u�3�����h��*�B�L�8��sL!���hh�o�������ݺ�_ʧ��.B����};(:M�w�g����<e�Ke�"g;虈��&��QM�`g	#�"���"�7�i(��{#-]��$W#��I�ׁ�~�)�#GC��n�C��@rSv�F|��s��ҁv�20_?8@���S�&��e����<[�*\qp����3
�E�ZNA�[��tE��a�������Ne�z<S�����t'�}���d'R��s`U�*5N�yp����A:�cx�k���_����J5��2�ҧ�Ґ&=�4�=e�m�N7ɮ<�/��L�0�H�����Җ�w���ys�73��t��S����/i��F}arl�����T���2P�J��QV:�Vk�j2{�|@X(�n'�8��i��R:�|���� ݢ�H�g:J�	{� �R.��C�"�Z��eD? Ȱy�?{�
�Xq��K��+���1tGG���r��c��ҟ,�S�}��_w4ݣ�f�������s-8���D&Q������xr˃S��J�2�)��n�?�	�5���N� z�)ԍ��#J{��C��W��E��A�9�с/4�7g��i8Q˕AB@�L;a�t.�pȹ����{B�Uv�4&��M�u��8k1���Xk�TI�b�<�&Һ?�� ��٩�;�~��&DX�~��Bv�.�������[���5��S�$3�M�Ty�=h��&��A	��/ /�#j�*.w�`��skNޗ;F��L���e�X���Kwa4�x�����`���8�|Sk�;f��w�b���O�)p���`n	��Tj|�.xOс���1o�L��pKA[Mj�B��oq��&7��XpL�[
�T.�Β���4V�N���G-�'W�׫��QFW�<�l��kG$<<;��b���I�
Z>���f�A�zV�������c�^�Lo>e��o��"��ǯ^o���PwO�4o��&�F� I����l�ѵ~9����.׶��5C���t��D��Q�K�2�@-��+`P
�e��JkV_\�0 -��dh#�H2.,�@T"��6��-���#�Ϡ�2��p7E���Z�n�4��2�:|e�/I�_�9�x^!9�_p4R�(]Ѵ�ډ�c�Ѣ
�"P�V7���j��ؿ��	�:���7}�\�oA���`�XX�Rn��+�Ğ_��d�/�-�o�G̥"@H��hi~q�4Ǯn�G����3)�SCq����(��%�Y���F��^�m��q88��x�z��s2g�'B�Di3��C��nDb���D�4��<�q�wЇ�J�!���A�����ѐ�i5�Z� ���nAW�����������/��D:޲��<�s��?����]�n~�4 �阓ɃEκ��:�3NhѪ��Iė�G)�I(d�4�ov{����g��t���z_)��o�;2
mCp��""z������o^�.]ȕ|��*<3�ן0�K]\��k*�oj�����\�L�y�^�X��[�	��>�C����ǰ ���E�C"d$]R��,�[MB8b0M����׶�����y�)ZTF�Xڋe΁0��Z2jp�B0���!7}ɡd%i���Gj�Uq
�P��ћ���B>�vuw܆F���s$�N��8��(�����s"�1����;d���Szb�n�͉Y�3��v'�_�b�9r���1�%�@�V �TK��&/�8�^�*��F�eCd���cr0kTU�%� љ=}���x���/�9$,a[A�B���C��c�=�^�'b� ,� Tvv�i�K����3���Y�C ��wn����Hs��s\Z�i�۟������U%��BHM[#Fǭɱ
��	&��i�m��9��H�ҍC����^��
�ݓ�c�8��W��h���ӑ�}&���w@]�F��>�%	�W�0�[G����\��*�	���2���哊�4$?FW�"�W��x�_�V��F��$0w6�
�.���A֙�#0����:ͮ�S��k��΂���ٜ�T����3���g�7��y���yb��D�p����]
�j���a7��7��#�Vyk�j=�
c2��!�h8�Č��6�`h[C6�/;��d��a�j��kA��=#7�!i�_!���g$)�N��]�̛
a�ei���$$Y&�%t/H��	;�j�|�X*��D�x���.���%��U��'���>�5�f�8�;m��y�z�^L'�����JߙY� EB�����[��F�2�z�^e�u�|��.'�&�$s9�>7�L0_,������ź1q����o�\�U��c�[�/@N��fJq~y���`��O⫛����i��1]Y����!�R(�,�;���wsP�2��u�^�#����i���ލ�x�������o�x(j-9�'��I�>�I��__#��c�A!j��
��]Ʈ���$z�7�1�nW�h��Ь�-:��jf-��UEWu�m#��0�S�/Bz��;J�sG����n+[^�x�7Vs|�W;ѺEȭS�;z�3<z�f��a�L�� Y�1el���SzF}�q'�owS�&�8����3U4/�0JL3��3�U�:��bA�V�OǢ�W�l~���M�cl���O�;��-�z�~}f��d7����������r��D��v����=ǳ��n���q��ސ����6Zn� ęo�o�/��=�e�c��,A���u����0&�"�2)��#W߻H��̽G��Hq>�kʍ�.�*ѱ� +���n`�&ņCkq>* ��B��8�L�(�(%�~+�ϳǝ����;tظ3��U�\(�pCy� �*�����*>)��P�����Y*�Xw%�g�:�&s�l[QK�x���}����R�-����ͥ)p�HIQ^2��u�:�����ǖsւ�co���?H�jN;��4���������������i6����cDcڭJ�r�h���ɳA�w�Y��9���=p~�y�UR�K���H��T���	I��i���z0����~=� ����IV���:S��K�JS�(�����l����w�M���x@�r�䍉b3��.�8���om��H��|�ih�Z�@n���V\���JVeṞ|�})n�q�+�O�z8b<�b���{a��k����g���S���14K"�'{:9l�k��k�ʡ�v�;��Y�Xs�Ts��77�Aԑ�O9~���(�� ,L@nc�6��f�ND��a,>!�z�����?`.�A!��S���i&f�x�}�rxH����W[#�u�=�2z���DV	�)2�4�գ�w���p��T�i���j�w^ь-��N�������MH�=���z�mn;����ľ#��Wk��i&���TGfi�w	�Fp�0����AB���\f�F'��G�i_L���r�JC4�3v֜RUq�J�j�p��/�D���a$������}��(%��XWY(�$�n������;�|`a�'�ek�r����
w���W<�NX�9�:��[TSu��]H��;)��v�O3Cx���޲wQ3&���1$:i�������c������9O+�`0HR�&�VI��茦J��b�t8w���?"�}ê�P��iB�m`�b�**O+_A݀���!��<W�=��n��2��������'x˥\�s�3�e�U�y���F��?׊�}����M�F�`����݄-A��T��'�����y��د��X��с��y��Ղ�p&������'�wځ�:�^'��� Io -�,��72V��u�7R�"j�0��dl��iH{���.����L���P4?¯��f}x����L�������8�ۅ�=2�B�����2�pà�m�ǹ����T=������j���<�NL��y�/ja��N[C�_������X�A�1r��@Bv|*�,�����2��w훋����?]�OD�ku�H���7���XRF��]��-!��7�5�Ƌz+I�c>��L�����y�|�I���� Ǟ�J\��`?�k'�T
,C>���0S�yB�2^鳽�@���[Gv���r'^wү��A�d���"{ϋ����+�z����[ߝ[���	-�Cq�����B���x�$#�3P��_.��)c�����ݽ�A;	�̎�y�kkq�!��iN�P&a
��g�����PP��UeQ���aF�����Ag}6j���^w?�c�u��"b�E�9�e�bvA��yeŀ���1�OE�e�#|�4�qbFP�m�n�<�C�^e������OV(�"�[垝��
T�ūr��pJ��Mj��������;MC�� ��r�����$v�~܎"��P�ao�r��ٵ�7�\����H��|��!��H�Lh��3g�|V��gr[��9��]�XZ���������i7���P�b50���S􊊿?1�*���nq��X�&n�e7qhv �O&�� ���kjzmow���m�P��6��Hq�xs�>����T ��D��<6�B�I^ƌu�x#P�x�l|�Y��E��S8Y�\��Y��ie�У�`>+jك{�����]q��O���g�~��7��\�$Z�c��k���:�T�1W��mg`�@Y O&�I���S/�MR����ru���3�dz
шY�j���6�}�f�śrR�HO�� �Z�޻��T���xH���{�ӏ�j��{�
|Q�̣�ʱJ �G)|T��� a�����z4e������A��"����ap}a{۩d�
K���Ec��֛�ʧb�,�x���	���̈tZ:�ΏMu������*�D�,9�Vt��&G=S1�m}1�7�Er�,O��i,�R�!���iO��t�`�V���r��,F��w�Ӆ�|�3aL-����#�L8��R|@e]	X)gHG�(�)7a@ܣ%U�l���/�3���tJO�g���fT���"��QF��`J�=�:	
�9�W��9c��iZ��ؙ���frD�c�K���*t���X-x�ʰodu��ZXn/���.�^8�w�$��,�{Qe�ŊvRe1�j��*���yE/��㘈L0F�����/}e��̨D�WF���-k*<� �3�\=ۈ��3:a����cQP��5q��N�?��H��ʟ:C-+������l,���6�	�	�Ճ���*>3ݖᛎ�<�z����0]A[ ����6*yږ����S�n��j�,��'7��� �g�x�t�C�;�Y ��Dc�{%�?b��A�xM�h���p���@�pQ%G��R����j+�j}Q���8.��б�d=՝�����ؾ24>�")#v���[�5�5�݈�ބЫ��>��tY~6$�ء ����F�wa�y����+Z�_�k�AV�z����$���@?���)=����{�p ���g�O�0�1�����Q	�M��:^��w�T]=;��
�tR����0W�B��-��x7G����-O@�)��k�����E[�J	���[d�����e�
fZ[V��]@�PxR(�<èꥨ�g��G|k�z�.�_�0Em�w��?�����)w�51�VE������vs��ЃLJ_��qR��Qt"����7v�:���c�C5�{p�^]=�BOԼ��v��\%�^Ot���j*�7;^]�6.����Gs�J��O�S��K��F���/H����il�ق��:4TB����~�~���8��Qy�0Y�ݜh�}^00��Q�y����nq��M#�u�Ā�����̑��[��G�;�d�f^�E@		x�s0q��p�漫�/Owd^��i�[���W0���(��\V�Q�����L��ލRRI��ݫEuOG!�|�3d�nӿ�^�TN\���̶�����2��Il?�.�9�{6������%yz�_9��8�[,.���T�|��*�7*<��e����q{�7p(G�ʴ�=\I�ir4h�Sb߹�l���6AX}���g�Oo��qλ$N�7���[��Rzf����Hb��je��䊁)��B�$Y�	�W� �}M_� l��>V���6pެ%�������H��(����.]?��,�PX�O�??6��!�"1o��\��چO�)��2�"3����'�Ԫ�pP٬o�s�D4-J�|�[�M\{n~~��K@��{.w��H���B1��֐�O�w��<�6�	3�xo��u�'2p .��^&F�0ՁR�X������ǰ������iV��m�~�Ȟ�i����-N�T��V�u%��1����B~�z T��i*l��~���k�$y'���JݾcQȲ�ВS�e&:6� ���D]Q���JF�BZl��)y�I�~�mtO��-@7Fx�_N���E�s��=���ʱ�q\�_\c�� ���H�c��+�6���x�u#��zh����n	D�dWhb[��A�v�0*�����	`�����b���o�Mw����z�pN�Cz��1I΃Ʌ%(�&���lz<�^��Z�o3WVXjT\�`���qn�V��Ga�ɬRL�܀��q.�%4��um�V���hݍ�\��ˢ����	[�;�e�>�F;˵�~�2�S:/�Y�WW;K��+�~cU���*Pԩ+k㜟R8���Kwc��C�@PJ",�*��~%R�/T ��G�8�J���h5&���\��gҮ����I紬?�־��Br�T����!����e�f�&�������Ij�m27!�2�N��~�nA�@z�T�d�ρΞ���Y^��R?p�=������3�y-�jš���FB�-����M㙏�YQ`���&��C��$ˢ8�߀7^����֘�����z���3��m��S�|���	�%�������bZy������d��=���72-�Ek���:������h7z">MB�Es5'س5Bͷ94fǤ@Z�6�$��,��w!���89���~�p���M��{tyȶ�m�sD�����ki�T6;:�{���75j���)�B�˙;ڵ��b]#�]{�P��y�u���wjY<�����2^,a/�X��gxbc>�D �|�wo�e���n��ط��wqo�/:(���[�~�0y��E�y����.���g&�/�DbU�F�ѯb�}���V��H��숄ͬ�Hv�n� �VGз�R�~M����d���G�d��V��ʩ������7��w��"��@�6�F��왙˩��AZ�@�7�c\�)��^�-��:3$C}7J܁��_}q����x��_��u�Q���#�U�X6�7Ir4z�� l����[��݈&A�n}���nc4�`Q?��|Ta3�9>�W�f@��E�4�5��*'h$b�P�zHː0Dh�Y�A_��[�#XQ�gy�,���%�vn���e��m^�&�&���'��n��'~� ���=ۖ$[}F�W�QH&��FM�-?ɕ���9ہ��Q��Ӌ`�<'Ŵ�N��ߕf�
�tvf��W��hCH��&=	��6��V�l��jE"r'���@���䵒%��7T��N듚��8g�Cqky�~X`��bPkI�3߇V��;��T}�.�\�Lɷ�
��>����֍|���f"e=ڻ��]iY��.��30q}�~b ����A�0S���_�.�(V}ޯ�4�kGn�[��U7���[[u�!y���$���$p,ы�-�m�I�5v�.��RZ�yD�f�B�͛�E�X�XE]�7H�a�M��d�!���<˵���p�������"��
v�����3�;���W��)$�t�>)u����E��õ�
�}�S���I�S��gPF��'7>(~e�Ha�R��-�S��5.���u��DÛ'����m|�E�J����ͣ�ō�&�#����t�.P�c�?��W���S*2��Bq��|�CA�z5�Z,��Z��^�?�����<} �<Pc*����Ar�B�����c~X1���Tb�9�L�{��ۆ ���8���<~'�җ۸-��D��=kAr�$�(��X]Lѭ��%͘����$�  �ƃ�ADq32��j� �ouS�+����M���t�.��� ��Do�^���w�B��R,�0����*�pv����4*m�}
W��x(ܖ��l�������d�N��n�;�	\�o�x��[XJ���S�M�$_Ԋ�Ӯ�%��J�,M�h�hڅ�/z��}��e��n��r�9�|�4, ���V"�˽���g��c�R�N�n�3�����c#jtpW	��Mq���F�ahd &:�x�]�Z=\��nҞF��l�}���G��q���~o�%�������gN���iY��L�ף�X�AW DzD��,��@��;�h@�0�K)T�1CY��zX�>���� RR���w���Ʊ�6V�̀ӹ�,nߡzE�xί"\rGk� �N��*2��ǘb�z�'�8>yfu�B>:��V.�b]�B���G��v6,CG�";a����7�Y)4rU��k_����bJ�L��d�ccSet�a��yC���3��[%PmYh_4� �\�)F9�*w��r�0&��DE�v�Lrݖɚ�'�ڇ��C_2R�*�,�\H!��[���h!on
��M��>pq�/Y���$Jt�X����\�7��v�Q������pw(�{�U��_��7?���5�w�P��9Rƻ�ay��jYnx��� 2B:u����9�Jk�D�o}��GCU�ȓ��0P�{
�t�ح���^b��p�oφ'&g�}G>�5����-���i����,=Q^Q�P�sr�	�˭@�s�|� �&M���Y�'�ݘ�G���M���$�|�(SS0٨:ϣ����+��Px����J oT�>�T��%�>�-�|t?!I�[jq�G�,e�H�zȽaE��j�x!$�ȪB��SK�u�������g��Ю*����~���1|&c�88�&:���PP�Q���#�Ս��z����d
���V�nf�jP�+?ӿTFOc-������m�3}��>�FK�Eߠ#5�e�k�b�K|m���J	H��h�A|>��qm�_�/�J����f��\�KL6�Ju�Ű��e�˹�A9�p��
&�P���q�P�"�Z�s�S�wdǢ�ɯ"�k�#�!��y'`Z�J��6�zX�{_\�H�x�K��*�ҷ\2��4�Ůe��<��	L�[M�_M%����}D�W�z��ק�)Z���e���f�	
��?#�^�:I���kf��6WT�*���hY���ع��� �tΌ��+3`��x�8� ��X<���Sb�na�Η\5�ʝa%X��7�o�&�d�7)Z�����lОK��S��p�ּ�����,�^��
�-�֢ 6�ae����D:��S�hU����H�Mg�w�ڜ i����x��Dq�����c?������,U<�Oސ�يD+"�Q7�m�&�̥9U�`A�H�x~� i���ћ!��:0}�kR�E*\����N�N��N���Pn���� ǉk�t����8�}���9Z8�\��9�z���L����^5/qORt�Σ<J��&&8�	a=w���̟*q��Ã�95�Mݐ�(Ab�w��`�?�[���b��I���������鉢۹�F��%}�X2!lf+��2�"�N�A.����[��{i���ȯ5&��C:�eP�9HD��7.?bw�K���k{P����\#Tb2>`P��H��&"�݇@�-��R>2��+7�"T5Ŏ��\$�ʦ�_��8�� ��8���*�Bϐ�!�RJ�/=zJ��Y�?�����$��2j�rS�"e%6��0���M���MnQٜ���"��7��[}ד�U"D��<A��튍CRo�n�؊�^&2_g#n���^knm�g��T�Np3����	�^O!x��܃�y�%�ӄ'Z��ӓ�9��*����r%�kM!֟���P8z�³�"9gb���`�no�	���U&�`p�y�e��5�J���t\��x�.�����B���
�4�XM�+3�@֜�߿��e[����w�O{Z7�eH�Q\`?�1KJn%HE ^PW�E٭�	nW�ųs�w�U�[��oZ-D{�����3pyR�+'ñIo��阄�g�� �Ъ��R��/��;�l0i~�)e�m~��7Z�[���5�W��^�+��M�(�P�Q��@&����i ���68H�(�[���ZúͲ?�JE����-Sgl��Ӄ3��+k�t	��Y�#K�a�
D��q��!�k�JY��v���9�*.B�D��P�n[�Z��\
�c��bC��f��x�O����	��{����t����b++0�4�r}�B|ٜ7��#�~l�h��&�LU��R���&��=g�	CǊ��պ�^�!�9m�Q��P,"�g��\w�c	�k&(�}��v�
���h�#��ч`	�-T21�z�o�r��_ I��� ��}Ӧ�v�f\�]=���"�Ŗҗ��ƿ���:q��9R$H��"�.=�ZZG#�[��,�oc@�t�L��d�P۰&���t�� U`��z,�B����o�x��o���=S��ߠ�����SaqDU�Z���V��Z��sB��eM
���D��uJ�0z��l�|q�&g�XZ5�wr!���ؒ�� E�8P��ܡ4��a�9�AW���è�7���Rw�_���UU�
����p��g\�=�R��A3��Q����Ar,�I�@{]Ԭ�I���j�vo��O��.1<�\����M���b�s��p�h�ea�E�n�
��,p��y
䌓�OJ=۬��L�h>0�k�0T10��n����'N�8���*~ǹ-��z!a���T�0	��ɇ��?����Z\�����/��q�=��2�H�m�llll��;��خw��Sꎶ'�J
@c,ՎC)�F��D�����3����->���I��ˬ%�)$��A�i-��s�W�Kd�v����Ƽ��z�d�?Ԇ
�7GE-��Qc�w���hm~0-[L7䴼���J{6���2�[�/��}$vd��د�,&B"��N�N��:}*�DB�������J���v�vPo��j�I,��Ap�>��vcX�f^9mN\9�^�P�yS����{�(�s��lג�)��n-M��٨yb�w/
�ޗ��]�������'�� @XgH����͒�2��Y�4�-��Z����,��~#�7%����E�p�A�YdT�	���OKz����O�G�+�����zpJ���ޛ���["+�9�)6Uk�Q���
�p`�}1�.����a�-��!hM�QW�c��B�IM�7�juH��8f�îQߢJ�f#������ߘϡ�
v ���:�q��pvb��I� ��d�!Ar��/�&^!�趴�/tJ��yM�P��G�H$:�G�Y\K�C�쮫�Z��LC�>iϴ��ȄJi��3F����{R������Nn=짌� ʟw�Q��j�)�:!;'���Ɩ��^����UEџ�5{4�K�\)�U�����l��*ax�P���F֢�y�5��Cf���;��C�Jd�p7�nvW���z����L�t�iN6����b�����m�ib�Gk�Ŝ�3y?�*ak�Kl��*ԍ|>�by;��;�XI�jN�]�y���S��W*7c�QK�+:"��g���%Dc�KC+���L">t���.U���ݣXu��N/���8n-��#���h4���T�"Ե�	��(B���Y�X;w|M�f��*F�8OF�\�|�F�.)> ?��S���f���/�_��|����~v��4(X�۰�7z,��݃*U�������F�R���Gh�h�����^M��'����[�#"��J��a�R��Z���m��C�/�,�w�ͬi�#�����:"m��[�X��R�6'/����C����H�"1}�K�o֢&�_��q����w;�<�tG��v�b��rdk�
\��9^�)k__' ���'��ڸ!-fF�Ki��m;J��^T���;�5$-@	7��m|R</�֋���6R��Wǰ�o�S�,�)S+�dX�h�Oi���s��"��� �jq׸qo���(�I�������"p��x�ז��,���v�*���07۹i��+����0��  .
	��gz#����L���|����
��6��7e�9�JO����1�:|.!��SR)8zϿv��H�}Lk���U�Y�4��Ѡ�IP��	h�6�
�|��7�M�D�̝Q�&r��W�r����Z@�7��U*.�6埍Ǵs�~!��&�d�92UX��!3�<`�+��z \��-�^Q�@�LN&��� P܀����U��)]O��y�;�q;/������d��|t\�~�wA�q���j�j�3���,	�A�%�~H9|X���# ������p9bP��9�B�X�H���xK�����?�I�Ġ�$����c&&�q�>� v
��X�6/Wc��P���^/��l=�.m{�)!;�dH��%܅'��BN[�LP},ĺ���PKg-W\,�?}��w��ªPiV8��/iG��ڙ�O�j����a���­��j����#ư���.�N~���,��o.ly6�!,��4�\:�q����7��X�-S��O�ou`�X�mN#�g�>�i��L�M��c�t���6��k��e��P22Y�������?�4���pY\�JKS������V=�GK,ˀ�bq�Ѧ��Ů/����f}���K���<f��w�<���WS�,^Hq)�Ȋ�O�-�<���o��Z�'�,B
��i8�<@��դ�/�yfW�����L�,sgL=o��?�./{�8��'�����b�����7�˱�����'�C�b_���g4.6�ƿO-�5 `k�1��1]�ʉ�j�v��MQ��Q_�2��FG�1yzϨ�3��̓����ǀ*Ӆ�����D�� �U�+�1D�D|���Hvni���ϐ~�
����Lg+]~Yz�OZ/r5G&���v��_�l|J�6~����l�i��!�P$��ӫqt�8�E1C��-����>��w���v%�0��a�Y��^��K����Y����t����0���D�p�pj��`�*�}�T��T�L��Y��!�_5�*��&�ul3��z<^�a���Ǘhp"(���I�Sn{\d�cX�~B��O������gw���th�\H� R�uDJ�곍��<����a�g�a�mxT����!gxl�Rc$�F���R�9Yo�T���<Z��Ƃ����*�Vɝ޴a��+�A��j��匟Z�9��������e�, y ��������j��݉%�[Ǿ���g���$b5��*�t��jX�o�6 # �u���¬��x���Ѣ �k��
�J~���Py�h�/���젰��np)~!�]�IQ������b�-�Y�7�brв��d��m�km��b,il�kI� ���O1�	%��<���p4��m�&��xX�L)"b��wA���h��$�\��[��z}�v�F��cM�Fk��bUl��!�k��"I���}>^�j��h�E�FT�.͘��:����ښ���pID���r�%�s@�����8��~��;����o�y���w�8j����N���$nw����B4D�������h�ֿ�u�9�*����
�[�?��cS�w9��|\9Ŝ@.� ���C��V�t�H ���O��ס�F�]ZJMǀ���f�2�6c�ӄ<��zp,���Ƚ��YN����(4t̃�+i9P��Ek^�jD��J�<��?2�R7`E���@Mg5=g�{���K��O[�/���e��TT��n{�H 9jR'AS������VR�L���$]?�a4)� �R�+�i�DJ��Q�TD�1��i��^`H#���K�f�DQ���&ͱ�X��s��l�a�����C��7�"��,�~3�}P������ۼ@����P \���[��2��f'�.��z�z�gk�̉l�[r6�?�8���x��w=qF_�����A��g� ���I�Z�ڟ���;�L��_�w�@��B��k��$��:�32����y�������߶9]�U����[=�C��2�瞚�J{� /2 ��i��-Ul:$��o�=���%��ʼ�˞���0��Y��=�u�F�/���o;VY�@n>�������CS�pR��*��AJژq�`��H�g�G�i�щ��o��(�|	D�AC=�Ⱥ�����k's�I]�ĭ�YL�X�t��9�XQ�8sx��X*��z0뱌�/G�O(��
������9�	��fU
ޝ�tm��,�2�g�|�<�[�զq���y��.�ǂ��O�X�3;u���'�y����:�'�h2G�F�!�H��&��|�a�+l�W����T�W��c�I�bN���G�3"r{~E����i�����u��i�A����aXvŃ�B��F�����B��rѽ�|�Q�<�lt����y�@��!b�%\�5�yLD�IO��#AaB-�˹c��o+j��dӋ>���
,8n�Ķ4'x�X�������y��]N��o���p	�|���8���m4o:��+�R�.U�Ӑ̟-L\��>�y����|�s�>���x���ޞ�秌��)m�?t�Z�a�aԑ��T�kG5[����\���R%ۇ��r��I��D=�!�8-�Lb�����"�Y�R�T�2�v�V���@�ێ�����9q��B�E�$�h$l��� \H�Mj�@��g	Ti�x��1h;�����"�{G0���SQ��2T�Z�a��[��L]���	 ����[AFסPD�N�V1�Y�̊�H�-A?�
��-=��*�h/�v�`��I�b�9�}��5˴���Ev�a~+M��,����H���D,}X"5�C��d+5l��d���Z��[FTY�&�־mWf�{��v�`����!��4�`�82�Ɲ6�&w�RYT^㲋
���8�U��T����s�f&n0;,�G��$�e���%G��ii�
��1m�b���_�/�*k���}P���5H=z��HU��.X`fM��v˽2!U�5%��F���p�ʽ�ٻ�1�j�:���,�ɥ1�Т��ŧ]�*�a�55]'�b��$�3�!ƆE�<;�L�
�5Y�+�{��{�1a�kKyd\C��
���a��Q�����RrvcL���F�5>d�����7�W�)[.j`{�u�:� ����^��N��[�����*T���t�y�Ev�����v����>��s�ӂ�Y[6���ʵ�}OX�]=�%��B�ߔ��a+mk���g�w ��na�o-P����v��yI=��°��t�;?r�N�q�
�~��J�@�{���t2ӿ�w�[\�w�y�G�_���<�Jr��PG�%��Y)�ϋ3���Qt���G�-+ͬZ��S�D݇s�VX�;^JP�a��vv���R+��{ߌChzʧ;�ѮFd	��w3���!���M|/dW#__���|(ПvbrrI��?o�`�B�0�h���R~�� j�	�����cJ�c����N�u��4[�y��d�P�,�ԗ�o7����»���yB=�\��� ��@A��x�}&m��:��h���}����x��]�_�d�:�A��b�^��.,��@u>�D��4�F�@�ۏ���"ə���/�4/���D� ߭�~YV<�,� �5����A{��I
)�q��-G��hs�bfa�r�A	�_���'0��/��>��n�Q�庐fc�ѴT��3�1�r}��SM|Q�$����g�G�39�W����
o�yR�+�J���I�̯�w�0{����⻚�n��\3�'~�ቑ�]z��\�|�ā�d���A��h����ɑy/!:$�n���8��=?��Tij�p�7�qc��iS�]hi[!���&_�bX���I>�^ـ��ȼ�rϱ�Sr�/��������.��R`��B�Ǽ�-o�,r�q��	:�x��-�R����3a���ü�O#����	���W��o#x���9t;0��q���>����"�$<����ز�ygwϊ�ܦ �����i���.��^	^���T������-�1�bۮ6�)F�����\a�[++�ݔ�@���c�0��J<���1}�ץSK1�T&�YH��۽�&#jp)�R@�2��z�t6�֑����=9�Bc����GY��a��Ȭ:������j�59��<�r,���ȸu�!��˚#��?���2�������q��N0HWl&��DolCUbĿ"m_�I�L��8ϧ��O3��&u�/�}��G�ߏ|Tv�yOv4(���W:�s"}�����7:�&��D����Tq�R�<��Q2����}���fR�SP�>������H-DwϩF
9o��	�ݛ(9��[[�Z�]�+Xc�weG��5���
L���4e*�P�<\���5`3�D�C�1q�w�`yN�\D�_o� L��4KWO� |���'�����HU�r�`qﮩh�!����V�T^F�N�hＶYϑ��3�C)��H�ω�a_��@�A�h��)��Ik�{�:j�W�:Ҹ��z3
&�	�y�0��������@W`�ͪ�g�;�0K��o� t�[o��l���T���BM��ww�M���P!dy^�cv��}|��88`���:��������.�k��|�f���B	����xæ�����7B��5"�V�v���M��5H���:Љ{J�l���!���П� +�1̾�x���4}:l��7x���A����A�k�L!�oM,i����?���:A���y��جt'D��n�\��M�],��7��&	zt��^��ǰa�m������Ia-E.��P�B��%��fh�{�F&��S�
�A2^� ��JB0<�`C�ġj���{í5�̲Y<B�����"i�Jپ r\^^��pu�Ea��	�M���f�(O̲�H�/K�\Kusm;�Ne�&�5�d-5� ��Ub���k����;=.�䖪��S��s�NlU��0��ZP܍�J6ӗK/-0 ���i�����c&�{hp	k�W
���6�ɪ5��>J�>�a�:"����RjdՐ�^D�zbY�+��~�vy�`Ɩo�i���H]�]~fy���;t+R�������?냤���*`�J��s[QW%��nE ��&C��K���$O���8��� ����
�n��+�!K���r��>��F�7:4t��^��լv�uC/j���cd݂�oV\R!�`�s��lޟ�����e9�t~�PsCW<NsĖ�6��H�m��+�%�����黜�L,u���X;3��ę����N�7, � ��n��f��3Y%�Թ��)v���y1�q⍢���+��1��>�0��I��)Mu�,��C��^�ɘ�����%����oYUfـ�c�b�05/�b�[������������<~ �yy9]q�ë�+F��S�W7�s.��`XJ~�dۛ��2�43AV��׫��M��M���&w�dU�pE�^������Qʝ�8��!�x2�.��/\(�]�-�.�� xSE��W�'��^<���|�r����O�c�|J3'����݈!���k����8��e���������P�s��X>��0oE����.J��@�)�p?⍠`\d�v�K*`���c��Qx½�	�i=��U�?K�K�8in8.ΐ��2��M�-�Ώ2S�&|�W���>��N(LI�؏���S��J���O���=�٦̳�4�����j�C�Z�������jv���
�W�P�Qs�x-G·��؜QD���l�u(�e�vh����F���ʱ��3S�[u�;��ت��D k��U��� g����p���Mz�g�~��CL9M��x�o6F0&���yF��^x6�h$��V:��Vm�ؓ��S�5w�̓�A[��3�p�*�s�)���������쪉6ß+�t��=ي�믅���2��KU)�(y�7)�;ob?xE\2�*'�$-��v���NZq3s������n+f��bj���<4g�8�@�p��&�MhP����a���ǳ����C0D�u޷A���$&��(�ƊKPE�S�C�7-kl��Ar�q�n�i��d�KÉ�ɗ�Á"��~�xmY���N�9?��%Fm���zO��g��_Q��X�q`�-���d���4)�T����F�Ԟܒ*	��O8�; ��]�S��$U��=�Kxbl�k�g�߉�b�34��16Y
�E��K�щ���D�=��F���)pb�D�j^jn�E�\�;��u������Ǝ6?>f"U�H���������d������t|B!�*����u���z���� q�*P�_��Ë����@ (+}S/�xll���K$�#�Y��l;�A!�9W��7�@�Pdm�ϛ0o�JԽf���o�"��Jg
M�?T� p���T!�&l#�Q'9�.������:a϶�ُ,ߔRhJ>���֮owV<	�����U7.���r��B{	$����pA��K�Ѹ;�X�]��ZN�����C��?� #X/�7i�>[�?jv�K��-�	ha��D�tڗ_��)��RBVy����1
b��,�#��ԟ:Ɋ-�3��z���-l&���������e���?�+3�~+过�db�^¾�.I���5��`����D
�c��ܫ�.-�պr��+��<p)�k�)]��an��7k���C�R��ּ��e��3�:�i�-g[�^15���C��c��	�� Q��I���ؠ���Z�lɷ�����g�� ,�۸�����a-@78Eg�8P�4�0YI�P�[6���{ᱜm�~(�2|a���:�2�$L�Na��Y�K#�����&%�D2"eC����3$I�(�~�\8ݛ�H9�#�x�<9ݤ�>����֣
�#`����&O&��Rق܁�Jۑ�W6�����`_���J~H?ډ�J:���*V��eɤ�œ�P��K;��p�a��DN��3�x�%H�f=���F~B����923���& $tq���y3s7[L��7n�-�AU�{A��R����/�7F^t"R�5������*��Oq<�N^�Б�,��[Y��.#"��T}~���߂l2�����̕=����9��\_h��/�y�É�	]�9�����.0"��u�d�<7�T.��d�Ӵ��)a��Eb�Q���⨝��8�}�UA�@�>����a��*/�.�;�B��ۢd�y2ؙ@�a�8�_�=F���q52��)B��dI
���@>�T��_f��G�Q��ߖV�������NA�t��٩��/m�Mb�q�����&|M�-:��S���Ш�>頔h��h08�	Z�ѥ���ݣJ� 9�,"K��zE@/��y���doő�q����74e�8��l�<EO��Ik嘀? ���OL�JK�����N,��GHl1��+R˸\�N� ��:9����B
<41���.6�8�)�����x^���N�
:M�|YGU���˺^[ ۾��i�L���3�V�ųR�}���zp���QE��ܼd��kxa:��4�N�������X���߹(ƕ�Q�e�Ɣ4�-i���!�G\��h���Jb��뵾0\�hq[B��HI��0�����ۏ�5��u8��G<{ۺ�m�iɱ�?ԉ�\ցa��&;��]AJN؅@҇�^|t�QPj�_'.D�!���F�3G V�,JG�P������F��nE�ѷl)�>e�O�7�h�'m��?-E���u�\4��jm���\��ßǍ�,{�,��A-�@	)[*d�C�TGHC�eQ9� ��n�8��|!��`�덉�� X���;�
w�P���Lf˫�Փ"Mx.%q���Z ��ے	���**��������*��T���M,��	�B��A �ވ���iY����btL�z[z�bAAZ,��~!�J%�م�Pq����E���s�>&�y[���Y!Y����̥{�q�����s	��4���E4z`�o�\Tƀ�s6��t5�}hT�))ܰ��D��t7̞"�qx�a���*�Ǻ����C9둻��w:��/.B$�V/�^͗�U��Y�X�d	˨ockO4@Ҥ�߃�}ߺ���k���;)=q�?��ґ��p	�oq$C*]��/;�#������o�ƶ����	�@V�z-k�ԡ���S}����4�~�S�Q�2�Nw�X�h�k%�n%���4��('���v��FO��u���m�hucQm��%��((���1	̓[_��� �"I뗫?y[4,`wf��p]VdU\�5���km<����"��8R�"i�0K�X9�'���W V�`��6j�uX�f6n��یK��!n�ޘ� �Jyt�$}��z�6�y\��"���/2����ih��{���rԑF�!]�26"�>O�'��p�0<��-�Y��C���S.b-'���Y�Fy��Ê`�ڋ�C�t0!�Ms�Eq������Y?(²h��,�X��Z �A?'����
"SwAV��,*�9�B��:-L�9j�)7I���rB1�hmzݿ�œ'��
f�P�cx��$y�	�+oT&·N�;������4VZ̢��7����iI�R�1�jQ��6x�i�ө��~�_���
ZE��f��[	&�_ft]�E�5җ�9�M�uR]C�RɫDn;����4$2l�s��B�[�{��U�ؠ=_5�e���]W��i��ɕ6�����(�p4�+QN�/Z��Z��}�E�'�x��@�}h�#�i
�vޅ+ף��\Wx'��ӕ�:���ߢQQ�-���~1�y�a#f=���q��
�ͣ+�&�Z9t��ۜ� ��Ӂ�kH�xY$	N�ȉ�e|��s	;o�Si�����A�fT�,�3�Ԥ<���[�hiq�(�4�G�j��RL9=��o��5�6O��^'Rq�#�ib3%]���Y1	ŀ���8W���BLh�c|:��gC�i���,�*�^aE��ۉ��q_�*�����^�',&�7�#�m	��3���Uy�,�W�w�	H�B(�a��[n��]��_�H[���Q)O��u�ܓG:e*�Fx�n�w�:�5L#`X>	��٨�z�>'���V������R�9
m�Mk �����)�P��ա��^�AO��O�~?�Q:�q-q���H>�Ϯ���"�&�Z-~��m..��_ez�d��1�t�����h���y�ܻr�h���qd���<�Ya̅ �K�ڼҡt:�<Шwj�$ϢK�Itl��A_��F$G�s�,�R��b3Ӏ������®{�{U����|b#05+�]yph����5"�GkOk~(�����<����l�y�ۜ��*���a(���M�Y���J.�L=��߽i����е*�� �Y	=mt�Z��=�#�>Z��
G| ��'ՠ5��B�{��K�wv
�1�Bw��]"dg�nm�h�N,�����B5�+Μ���)��������O�|����xG0�n�
I��g 49�v��g$��dyG)����J���{gW�䶎L��c9|`�."�rz"�����S�}��d�<�Hl���[W�kZWfT�����p��g�/H���3��2����"#�}����v��4:����f��h���!2~�4V��p���r���k3�i���U *k	��' /D`�d���Ԫx7q���Hdc}gg�E�<܈VD:񖄉.�Y���|Q��n���Z�|AZa�0���?��S�!����GdA��ؖQ5��i㞞����)�a;�P���ݤv�0�ZI��(�L"�JW~8T���K��r��;��(���y�̫/�w��F����ᤈD�+ �QL��	��_W|�Y����T� (7�/h6x�S����-$�^��I���`(h�*�\r�|�s�UrUؓ��ku�PKZ�	�û��մXʚ^6���,���U���9�Xv!�+#d`^wߝ)�C���y7Q�l�:��>���B��~"������U��sS�z���j���l#sgRb<��i��d{;�i�w�7��������$G�So���4������f5������H�2�9.��<R|���ؔ��G&`��ө�0��#EH�#%�d\����}�ʊ��\h����Y��T�4܍ܹʗ`5�����|�΋��9w`�˜-�R�3��!`�c1����ߋ�i3�}�H��	o�:�Z��9xC���1�Y�#'{�[�~����	1z2�;���|Q&�v��r7iO� xDQ�B'!��/��pʷ���6Ԅ��O�:� �ui�����T�yi��:u�Yۥ}�S�}|�|_�E���E��HNZ9�t�+�IT_�J�hd�P���uᩖ�5*���K��Lqfk���@�0�\D� ��L���2t}1��;��w����U������X|����Mz}*-8��nwV�%,D���]�!�f㫚���k�Q�9�U��!��w�G��z�X�.W`1�F�T�`���yTm�]n����$oʀs����Y���?OB��^��%�o2"Aћ\�$*��5�{������Ѣ3� Fi���m3ؚ��In<�b�5wvMM`E�D���A8L���ƹ���eX>��ol�<o���1QUr9g�fۖ��W�l�!�8u=�	��Ua�M^�"��ۣ�F���������ߞ�0�;o\hy*�fL���]�X�%�"\��F�V ��w��͢ͽ�4!�옄y���9]�m�[���4=�Lȓ�ƽh�B��[w��dc��-%�@F͟t1k��Fs�i	�ޗ/�Ɖ���ڛ�ae�N��tZEk,Xk�%.�w�p�%+݆�A��ICʙ�uc�3�~~$�M;B�����4�p�����"2�3����H�B��ϴ�����yg�K�܆\U�GO:����,���#O��\Kh�*�\ΐO��@ɍ6��9�Ӆ�!�m�������.��"\�.�N�0(�f�3zVel��{3�)��7����a���r�_ A������2`)�=�M]�A.�sg*7�`��L�0�A+7O���Å�x�! e��{��n�@�T�f�x��1\G���Q>KO����B2h�����	.��P8�?��6�;\9?�vQ褊/�L�S��4��W+����rlo��d`}a��2ۮ���?,�\Y���!@r"����U��rƼ�e����~v�����h�@P3����)�@�:e� �1�����s�~�_t�c $�y��[�Q�sd��Jlj��M�g���"�23=�Wg���}G#p��ۧ`/�A��=��&(�:�@$��h1�3ou��O	9�a�;��ebRX#F:�w��N��3JY���K'c��pvv�`���J�4"LZSB�i������5��$a�R|�$��m��`��\`Y���3���ż��H�9T�ߩ%��&��$�)���(�t��U�a���x�RP���lo�4y��Ǽ��+���Em_j��c�?O1��.�x�u�06���1�Q�S���Y��.�^TӢA�m/@j4-�ta�$5l��[���7cl���s�#��9��)�ݰ*���}�����3Ǎ ��%�Lׇ ��i��,��7������G�:��+�Z��F�8^�ш� 	1��$�z~6�g��g�n��&z���`�a���w����C����	�m=����J"C
�ĭ�ދt$�����1�)a�v��W��M���67��T's.��j�GQl<��0f,0��Ŝ�ٷ��>��()�`^��|)�ͧ�\�oG����{��򻢮PD
yg��t6]� Z*Bf��.%g�\���;ٲ�u#�$Y�󬰲�b%�7R��^	o����}����ۮ4�������?˰�v�gQ ��iX&m��m/1����3�r5�=dz|�On�Z�{:D����*�DAI�mq�8�q�s��A�j���3ɲ��]o����t��sc��W�/�R�h�8�+�-�y�6π�?�i�{��$E��2~�AH�d�Q��3f"��At�S�L�Isk�]8.����E��5�I�9�N�<��&���Ҕ(	Ɋ���?L��������TVO�h���	F%�C��
�zĠk�i��(��7u� ��m�3.�p:ʰ�y���V��U�$z�!8+�E�c��4`���Va�`�<�2���lF���fn�k�a���!�OE��Д�Ձ(w�#���ܑ�h��
��Jf�c�^�f����~�J J��E2;���_$+�%8d��T��>��R~=�n
�K���"��?�Ai�Hr���7ڽ���NNT"No�v&0|ʊ��#�K�|o�C����V���E��݄�18K��9["%��C������?�U�	*c0o�5��D��3�\����c���m�͉�^������o�2��Q�x�c��-&�.��5y6FT���3�	
�x�4G�P�n��2"Z7�1����g#���i"n��3w�����G.B� �1o6�{V����ǁ&N�B�( U�Rp!k�Y�4��\�����k�#"����^��3~ �זkS}{	�&�<Z�6�X����A��^&<�X�N��3ǃ6�K�-,��%*f���@�����!�4����c�;��GeA]��hG�"�Z!	��޹h�W7Zf�Y��U�v�p���>�?�O�牤@��2=Ē:4��'�Ao	6���c��⦃��Ŏ}_��#���݌0Wy*���:$����yk����>�����7�t�5�+�H�;�v3\fe�>v��'�d�lG��T�'(:�I�D{�Z��~��KŚ�^�����'=����ڐ?�Q'�b�kan
�0� ��%"�B���`��2�%�x�(���/B�Ϲ�v�P졯����T&�C����c����<xWF� Mv��� :��Du�l��t�t�pQ��Ϊ'���G�5�6�x?�<��8��}�02�&p��ν�E!԰��9����a����p}AOv���B��)���^���"wl���&e*b��_�.��|9˚�� KT�����Ş�ĥ�E�ލ�`���~���R�9T�_¥��Y��,F(ᶕ7�1G�yN���44�� @�E<�U���3�-�׊ͯ��zo�N~�?�*�P���g�.��>.��~|Χ�t|�Z�}������]ɲߘKf�v�m�@dC�*'�UͿ�Ӥ:j��;��f��@���2`L��������$��L8v̠��K���xGP�|e�{sU���.��M�@��+j$�2^��D�Lm�%+WO�K
�v�K���ϙ���p�Koh�RJ�}����I�H���
ḃBÂD��9�?HDoI�#�f|>��k���V"�Ⰺ��6w�\6cMF��J�)Ԗ�0�X�&���tY���q%7�u���g�cM�}`����SϢ�'2���Z�.d.�e�]�O��R������eV��&�f��r���h
*��ӏ�܉����6T�n|�T0`$�]M���=�l�P�|\��م ��M����3����0��N(]$v���7�7�v_�����̃�H�dZ.��&��?�C������� ޕ�'�aҐ��|��*SV��>.���{U4 {���j�G�~%�x��,��W)KX�K�6�׎��-��mD�K���[��*ו^�0��l��p��rޡڕ�tө�3���%�>�W^RG2�4�:� �.
�hYJQ7�fC^���h��|�DqR=G��R8,�,�y�A�QR���1s����6�x��f�� �����3���9�A�es����;/<�(])���ܕ���K���:��g] �)��N!��p�a���k$f�mH���4�q����]T�ϑmΧ|�=�@r�CHG����^K�{W��G�ǓԞc��]�jE��3uM��NC��H�~)����y�O:��ē7l��O�N(U��hcڳ���5�S�M|WZ�fcHk�?����xi�ϊO���#ƨ��1����ˏ�G "C:����)�q}y.�x'.���1��5ݩ��Z��ڿ���ot�46rd����*���W��kKh�dU��,�>4-%�>��GFt�_4��6��א��[�A= E��d�oj�&m����	#�O�;��l�h�P;]�/`l�ν�q!*��m�����4�?D�S������b���@�пg�`��U\�-�J�I�������D�-T�rqO·�t��B�4����D��1�Y�˔}@���&U,A����tҹ�U�����a�ߧA&�[�U��`��Ѐ�w�8�ĳ�-�+	E����%�LH>^�ؚƈ�C���p
�~M5���j��@{��,-)�AP7w(���5�\�O����>.�	v�P�Τ���1�3?ҵ��,;�&�NP"�.n����<�Š�F(Z�J~8iX����&�)9X�ͭ�T�m�I�*?&ź�zq@�8�e��$g��#�f8��1X�ǧ��5�����̖��E�f��&�郕q*����������6�qn�������d�c��|�d5�}���R�]".�7B��~��<X��P�,�Mؤ�յ���f�7��!�eHV�(�=&��X�8�y�\f�+J��O�g,�D�R{LN뼌��O���4'9���vX�t^�7�	�w����o�\� #�H}�l�	K��Y�D�a�\U��_����^���o�c���k9S7ۚx�� _�_��wy��c�_ݿ`�	��@ј]�L�ă���f�xS�y��~+�-?h���J����p�%/��{9�����k@j 8�	�o^N:W�,`,"9����\�����KS�0Q�od�S_m��������?��g��*>���%"�93,{R!m�D��m��Z��
��p��� ���X8���(݉���G��*�i,��vO"���h?�نNA��h����냡#��f�7b��[�������ɳ��B���DU��v�I;{._��Nh1!��'����.K`K�
C��X�H�`���zT�ع%m���٨I�5�%��o��m���pj�;�6�Od�9��W5�ԄC�d:-���'_8AB�Z��`QR�6�D���sk8���f����>�+�[�9�v�;`��M	r�U�s��t0��ߐ̺qs�ە~\A�}��@I�'J�� ���h����Ɋ��!�=7�u:��T���Ro���D�sV���B(|��
6'�Aԋ�ӱ"�Jm�i:��1e��' �U��h��Z�qT\EE~�#X�L#��l�3k5;y�<�Ӫ�?
+����)�b> �0�t�y<Bj���T��(&�}l�&�9��iULo �q1�D��ml(Q����i�%6ݠ�_�(pz�h��gS�����e �ĸ5�����^/��=�u�ـ����W	�� ���H�p���	��<<�8�x��q�)��D���8�[I+��M䗛��Q'��8\ȱk�����~Ԩ����}�"0VAs��؄��	���aω.��h�9
T{
׹?*�Ӏ���� �=|V���ڻ�2w��0�~(懚�jo�)�T�~�]�o�5�w��h�'�-X��B�9�����٬`f=��@��tZ��FR�f��x�CNO��X僇%*%xhaʢ���߀AT�7~�;��x�*��IIYPX�4����N�����̓T�b̳^̍k��7����meс�䰰󭽑Qꮍa���b>b�}-|%�A��Ar������[�yV_Q�8֭�/�+�07�M�����t�"��!��2ۮ(cзF�'+��v_y#e	��?")8������������`c�*H/Y�3؅�j��+G4@��xOϘ3�.�؏��Q4ߢ��"`�a���+�����k((��m8G=yC��sԶ"�ϣ�H;+���n3�8�-�A���Y(�T�)E^�-T7�\%���Z�@�U/r��1ͥ�](��=xv�"��qI�Lw�a��qʟ��%@��?��F�"�1UA�i^VA��xq��B=H�<�C��t���1����b�j��M��~���(:��+��^10��N򭈼Lo'�^Tq���vm0��s6+E��������^ZMX:v��ܜ�1#��,�f�CP�����ƙJ��,��>����y�!4�5��:�V.����]gH��r��G`���ڭS�8��S1��w�sBsXd�6�R��fH��V&��A��X��C(z��܈��ç�6#W�Vľ�C�=�!���R�\f�CG:6�����-��2X�M�^�(y(�Dv"殠����:��$
صo1��,�/���;p�)���	O%��$���8X]:�݆�ܓd:"6��bL���.�X��1��푋��
3�M��2�:naщ�j���Ө&��䖛1���O�P ���5��@�p��:⿟���Oe&��\�d���U�Y'P��l������7D�~H
��PFt4̠���,'�AQ�RM�w���tZ\]��R9��=���l�9���`vTfs�`�`,�㓹l��r��'͔�I���瓓�X��&��G,��5`�\1��s� �ئȲ��BDL��s�ӝ�!/�o���$6��,�?��@t��77
%�	n"!Jsi�М^ă�@��+n�"��y3a���S� "x�踄<v�?��5	u|��Lkۋn���p���^���C�ZRN*P�%Z:n��苪���Y0��_S�g���`����	���KJ�FZC��~s�(b�&�����2������Z�tf�8����g�E����� �a˜ ����Q|�x�x�F�{@��t�M�}ZB2�g]���CR���i)ia�cD޷U9��Ψ=�vD��(�wOuh��J	��5\e�
	��
�wS1�?������x�C��\zm?����0^��^�\��ӫ�@����T�R������B�
��X�_+�|�����i�_�RG���؞�����K�g���S����� j�U��a�������d%�b���7#�S�W���6
��_��J��2(�O��7�p!���E((cP��I�����O�K'Lbb�&��wb�B�$����R���0"C�L�?��۹4
���q�\&��dzs��)�R��ţ�=��`���P%x�}u���^���/e��`�m��6�<;$=��-��z�G�/ɚ+���jXmx����qsMqJ]{eE�Ue�/��-�$�c�6M�����VB���_�+��C����Λ�7e۱����cR��,�¯�3mY1Q�#ۣ;Y�.XgJ�����_z����r�J�T�H���]'�Deb!�T$�W���D鸙����LxG����HO���<�L�q&#��::�2 �Z:��!�l�-�}9Gg@K�u�]�c���y�ր�LC57r��	�[��l44�;��VI�m�׈���7hז;ݓ/��pz�����T[���$f6޳���ho��<Y�����0(��I(X�v�I�BL�ʥ=u�+v���Z)n�?D����T9rC?&�c�"b��,�R3����3�}Ӎ9��v��7V�B��W�^��b��������+�Im��^�/*~�U����i/g\i�kB���}:�*�RX|a��T*��.V�,�Za1�{�����|��/�̽O ����c�C ��/&g����GU,��o�4"VA&Q�s|·Q�$O7.~p.��嵰�rP�.ٿ����Y �`3���_G:�B��/*g�&E9�����hu�.!�p+0V��ry��9ϨT��/����k2���Uf��(�3���w$.��qB<!F�n~p�	��La���Fn��^�����W$���*�����5�Q�Y����5 ��,��m�>>]�C@�ʐ��i\F��b�	��zZ�i��q��;\�,�/��/��)$9y��P�k��b{�?��+v���А�H���\I���.ZXQ0�^8Ab����^�4�|d\�ϒd}*��t#憴M�{��Ε����~HB`"`ff�෌&%�����ٔ����Er��^Ս����Y.#��p|���x%�K9�m�s�2F6W��f��jҊ��#���z�jܡ�z!ubS�6],f۩%�f��n��9_��ٲ�\��������Xѽ�ls��7_3�!?�n�J�V&m�g�Z�F�B�o#�zdh�*�{+�л��y�TUb�*�,ʻF(�CP�Ҍ��:Ut00]�R�do��VE�"R+��)E����}��A�����T�~Bߐ�=�8J�	�vU�yL�շ��/�D�zJǬ��Sm�֫)�-Q�x�&���t��^��WK���Z%OFW{����5��lSe�w��M����#�[�?�7�%�H��Ԫ�Bu{~�1#?�W�FZ��~l�\��	���p��/�)/JW�I�b���NjR��7��V���0?�����ξ�KI��6�s�LP1��@3�2�$4���N9>/Y�x8ap��,���/����r����YJ�����TȦ���?������"!�����ɼ��[���$����~� ��q���-.rwݶs3j�L����T�c"3��>4���j� 'τ��I�+MT���3�]�����mb1%|o0��7�:��m�������=���@LW��	I�Ig�&��hʴXr/��&�������m�'jE��J=��qJ�G��x�Q$ck�|�o��M��l
���_ϰ�}"R�"~���������޵�&����6���$���V�ؐ��=�و�a���y-ѐa�)���%��k���?�'9|bX��9ӣb�,R�+�����|VIV��7�	F�W]{"_�C�0�Sq�p>�����y~�8${`go�/�6q������ڟ��%h(}�A�.��!�:D�`H0�\��K?�}�;��B�õ��&�x�w�oņ&C��M�;u�if��IQR�@%�n}�d�P/v�>���V%����1I��PJ!*po�
w8��f�V\~��J�Q��'��@l�4\����2	 `��{�+�t�v���m{�O�-K��D�_F�?!$Ghy��9��φ���/��N��ǲ3wSn�Y����\�'�˷@c�n/�~�����l��DZ����(�ǘ�^\@>��X
_�QV�L�f:�?%����o�Eú����H*�_ٸ�p`ƿp�O,��@N|��w'u5�����;���=.>��jש�wbU��ۨ�0��eW܉b�=8IJ��޶���[ׇ���פ�����&�
�`��/���tr����R�:U�.��gsmn��<����� �V�	yS�o2��f� ��R��Jc��
~P 8lD�������M����?ϭ�J��d�?sM�B^7��X�H[��ЇSe��}3iE�@�{�\#s�j���.޷uX魐�R۵��ԉd�?@7�����X �^�T�����G�e�Z�Yz�X-���i�|ʞC�(�Kfd;�:$� �ir�z������/2��H�S���[��0���q@�)��C�*:>��m�J��)��:�'��,]�������z�͸��[p��d%T����ׂ/�PL��%�T1޶eG�N�
cW6��5HpE�b�I_�������?�����ll�H��_�;9@�I��D�������-F�8��( �=��z+��ue����$�d#_=���,��
ĿbI9��{��4ȫ_@~��`u'Ƌ�� C�=⯢HW/��R�����2�2@�ZHI�ut|v?�4�_����/����/��Ic�˲^�t��6�A3�y��;v���$����\�ZZ�P/�R�{��.o����AՂ*}ŀ�2v)�$�n�M[�΂��C�
ǸcuEEX��D����?=�;��m̵��:�\֞�ىc�
��pd�_X�!	�ęm]�w��" ���Au��g���bm��"+��u�G!�Pa�7�m
}m�H:����W:�F���*�F���UM#Ї��`����������!1'�E��]A�AgF��S���%#q�oS�)�0��a�~��y��u��X�$��RPo�kMm�S�e�sI�	��\���|������,/��Ե��l,'�{�	
����������[�(��t]t�Oٖ��v�4���T"ISW�)c*� `>2��v�q�ΆNAݹݟŶ��'�t]hP�6���m�~b����?|�s��t-��<3�OI^��.١�C'�Z�|�x�ٙ�H�����Dd���l����WҮM͠ڣ�Š;q�Z�!]�D �;)t�M����m ���uã���Y�s�=�7cK��z��Wvu�M�ayY=96v0v;�ϊ=T=���hvý}�G��ʔn����W��5�E|0z�io�s�Z�`SR0��7^G��'�|��%�@�[祍OR�����ўI�,�4R-��׮���^'0J$�Ԙ��$�	|%��������rD�6��[i��ֵ��f1�Vl%9V��'8D��Jɒި��|�?�L����ޖ>t��z3ig_��Mٕ�yQ�����-�% S���ꊣ��1L��ƙ\��US����5k/��������U3��C��lK�b�p�Q<�ny������s$�[�#F^�K�a�q����A>�M�Kp_��QӖ���Ϥ��薧)�v�3�z"P�-�H�
^�|�>��ן��?�j+ߏ�K��mx�v�@�׫z���s���=o�bI3{w�a[G0z%�>b]�.�:9(���P��H\қg2J>O�r?��`��sxKA�<��%�伻�[������ƩO��8���鸱蓔���V<:�k�L�Sj�8��3]wUu� W<9l�I}�z����6n���sYx ߲�������68��
\~���#s�/����>0�)���j�ޔ�"W����}�F����YҬ��fS�/X[�+l�I�R��Z���'���g��r�č����#����v0�[X;4k�쭶N�b��ph�k��`U�ć�W�����*��J�М��zl�
�O�����/Vb�٪�zCh	��XdT��.����.{��vס��f�d��͖S������~:��$�ԩ��/��ق��RM�
�4 f؃q���He���'��D�+(���B�HiU�7��P	��|��+�6��R"��{:pې5��9Z���PB�&0ǡ<F2���$�3'�:��=G�c�� vü^YT�E6���a�w�@Ex�:�`�m�qRXԐ���|�X���|"�j΀+�7й�x5���[蔜�(�Mr+�'��|����7}/�z��a��4�K�\�����u]��0��9h�i���9\$$/���j������kO����FG��Ê`r����@ǐ��;�u.��7�\�t�A�N��cϬ5�.D���W]��+~-�BJ��p��a=v�B^�A���Mhx-�;�\"ѮT������^a���(�0�fq)�M^�LI	�+�lQ������|��X� ��-�=>�s&�-A�5�ǮTΐ�-��O��桗|��?l?�����f�t�[ ��<�J��������&�0�(�7H���T�l�8�}��[��f:.?r�P�-�2��yY2�o��UB��\_Q BM���k�#����
h��C�+^�f� )�9!�p'X��ˆ4A��;�q�?tX^c��F��O�jX��qi�����Щ�Jy�^���G��
��ǂ��J��"�=	��fa��C�q�	̓P`p���7�E�F^�~��|��ߑzf��������#�(y����QB�L�8a���3��,�2Z�k&�s�5m��N�ˑ�W�t���0����*PE�tl �:���"�-�Ҳ�V�O���s�l����և����h��1��;��Ȼg��PJo��q�����O�w�����̀�%zJ�vT9��n����h��%n�o��|�G#(3VI&mq����Ы��ɋo���U�*<Y����!f����V{{��,��J[��z�2ETY�LP�������) �J�m�U�=-ccRE�������E���K�2�0M�~���~��;��xt���=a9�m��P�U�e�c���_)���Ys=�_�rE��l�=���}��|�?�M��T��X�?�����G���O����}��V��38i��;9L��1����ѹ����#�u�ߓUq��@���X������vέ"���פ6�3��xqu�R�{��Z��S��G�}AD�r5ETx�><rν5n��+�Jsp��	~��Ν&mo�f���b':���5�"zN�a!���'IV���+y���a�O䠅��2!�Rl������>٢�~�;��w��+?�,��X��g�g�!{|9��1Ö@���Q��N�Ь@λ<�~���k�9O�
|�Yn�'4���<\m�Ϡ��l*�#7����}B\A������J<Bj��1���A�q�qȄDz�2�h��l�����C�";��q�bf@�|�Dh޻����p�M�L�J_�42�q����<�O V���2S�N,�2� $���,��[H�Gz������D^|���d��v{�30Z�%��*����<ǐ!�qܺJ���k'J̫�M�/c~�Y��w.O�rX_�?��?YVىcr�Q�y�Uuјc2�S���2�h��^ݽ�b �������qb�(��O�e�v����
��ڷ'�4�3߉��ZfƉ�%��yn�����sdH:��G��#�a��jB��"�VY(�W�1�IŦ�,X�JqO�B�a~�$~E�[tF"z_8�o�Ł���&E�����tҒ?P��5⿰C�>L��x����>�:\o�c8�Ű�|��E�b����1cc-9��!�*��$&����53��w��߹*W����Fr�q�K!�"��W�8�d����h�/���,$��Ӊ]l;i}�@֚Ij*�Q�������깱�Z��A��۵�����X�h��o��r�E�3�2SZ�wZ�ZG�շ�@�0�M���r+�8���(7Y2^Xn������v�d�Aދ"h�i�|a	�@�Ƨt��>�ٕԫf�����8�2�yWZ`�7a:�r��Ԇ��h���5na� �#I�Ӿ\�أ_�`#SQI�/,eTq<3��@zT6��`z{�r����?�O�]�hnm���Rn2�*b�'V`�io�OZ�=d��.��~��L�_X(����k9��	4q�h{'��i"�PN��ƄC�ZW8|i
�q�&l�� ��|:xRIE��Y�������/X�+�Q�+�݁�ƾz6��&��ߚ�S':�	��q��5g�Y�S\>�vP}�tճ�CA���a၃�b���f4�p�S/c�P���Ex�$x�]�������h��:��ki�?� ���
20K�?F��jʂ`�rK���X�������2�:#��"� �]M��$_sV}}ծ]ZV�Q
ޚp���4C�vA
���� �g4~ o�Edt@�G+4�K)�:���;ܩz�9�\��j�����.�#�l2��>K�3��A���;�in����!�u��)�N ���B4м��GI/7CI��~U��KGA^�n��Y�Dh\�?h=2�.�V�dWO�1
���Ci�G�<�t�a�y�@c�):�E��hR9�`2�w*Y�}�E�8<�,F��!�Ոv�ժ*����SI�v���]��C��'�20�(�5>9`�7�Jr1H�?�YZ�S�V�FFR���y��tF��@���J��!��"���[0U�C�H�4��:+n~�}u�x-餸�m(���s�� c{��! bH�3������;��v��o�/w��7A$�d�
�1C�H=�]�h������)4�V7X��͛���'ºSt���_#ܖ�����
;�([��Y[�'�n�5&8� G�& �O<A]J?^��D��
���pY��Х��1]��˸\�N}�L�4���2,��6���}iR*V�(����W�S�o���wа�^�8x���<8L���~4�$�
N���d���3��
�疑H�#�����asp�|E1�3�s90�%��vTIF�A�	xś�ջ]|�kO
=��Sl�k�"��	!.�S@ɒ��J�GPD-�T��'"���O���r��=P��r�#�a���p
c!����``1V��\a����B�,�����ך}���$ǼP�HI���Q0���]�đ�fO��p1k��F��l���	�J��Ἐ���$�K>L����6U&G��l7�_.E\��r:��~l� S���M����y26��ؖy��v=�5�܊��e�����o@DJ̗��}��F�90�4�Ռ9z�3>���:���� �$�4�4�܏pP���)J������ _�i��yw���Ѹ���Lt�y �� ���kԊ�\ߔ4�?�
�D����Z���������ƃZ���vD��pwjԨ�܉���l��j Anf�.�L7����kF��5�,//��e#�	0���:�D��ʈ����Î:d��:L�i3Y��̢�X�FW��S�.l�[�H�lG���O������G�3�� �犫%3�쀨���4��cb�w-CH��ζA"�.��� "�3�4ʩ3t�sN����[�_)�s
Ꮰ�ЖoTx�&���F���P+�)8�h%5ck��贁�Yp���ٹ@!>04���!�$���|�t���?��(�D|�\��uh��{;T>{MK���Q�Fsz��U����W.�صǠt�a��1���tƳO>!Ԧ�rƫ�ţ��ܗ�M�Tz���%]�s�D�]{V�Ke�/߽�ڶ@g�U�Z�7����\��Ţ�ո���x���;�+��K#�/F�e�ݬ�B3	�F����w��{��ɱ���&R��I��b!ⵝ���c�Zr�Uo2�:��i!H�1s�d��M��.������M������DQ�����W��^���������;�"�&��o�5�R�BйZ����xo�`����"e�rT�{3�xd��0ϡ��$k��a�$�? T|, �ִ�dῤ��0Qyk��r�Gĸ~�����[����.�w%�9T[�C�j]2��1��K���eEǟN|���أZ),�_k�+r�DP���p��.4��/6�^/M�땆Iy���38lb�ca��]�Nt�dj��A�Ѭ/�$�)��hK��N`=)�'*T���� 4w��s�د) ��@� ğ�JS�?��R���]�^̄R���x#�n�Fe�X�
p	���Y��"hi���9��+񝕣Cݯ�Q�z^����1�@ɱ�P� U0���h�3��m�}yx/�V�`���]a��D|��Qe�������`i���D�Ds�h<8!�4����:�����MG"a{�~�xJ0B��o֩�D[mVfLj�Jcݱi�R�er��6'�n���W;�쯕�{��M��&��K�تd����4]���½�B޹h����7/���z���h�EeBߣ9v
$ե���
����m��x�E|��b����E��1�y6�����	<�ʚ��y�l�����G�O[��=j��_�*�K��1�����)�O���Ys��^����Z��g@Ps#|�O~G��� <	o�I�%��Y�jU`�PbU)� �~fm��e�@�-�;��r�P�τ���?w\�ݗv�`ds��)�Uk�X�Ѡ�����qVUH�;hO?t��i��>��詘|,�Ý�!薯r�>���uD)s�	�i��W�ӓ�o���G
���M����gV/��
�]�#��z����!���s�T�C<��s�:��)"���\y��i�� a|C�!��S���k���3ؿ���dy�����;������wF��$��Ԟ�����꫃R�F(��C�r7UĘ�짮b_�ؿpV=~��/J֐N��E�Y6��E��Uqd"{\nX�b����dbZ�(�r��Eۿ��!��&K��	,�?�.F6-ċ��ܜMQO9�o�U��ZQ�
�� �u\����ܬ�K��z,��èƚ�X�+I�zd��>���!4���w����X���M�����o��JB��?��|�}�E�0����eX���#Mj��ЕD����8M�
Jg���>�K����.�����C��~�m�q�7���g8=�Y^	 ���/�(^�;�t���I�p|Q���+u'�R+�Y�w�5I�����N)�9�PS�1,��oY�g=���흨��&�>i~%f��h/������(e<@P��,����v6)��% ǡ?t����ہ�ϳ�p´B�W4���£V���
ޠ�l��Y#p�>�Wm0���Ϙ�i��g}aK���/�j}>7�!�`Q-,�S����>U�#8��q�tڡU%�Mi�����Z��E!+p��m��$c�%����ڏ�
���ְ����iы��9Pp�𨘚��w��qu 4D���S�㦝�����Q� ���O!����<�j��i[b��g(UjM2��2��ƟvQ&*E��t����$3�V�?��k�^���\s����(i
/�F;�_���.����Nv~xq�;-�OI+�tWcB�Z>b;�<����e�?ԪXg���7�/��Nd^�m��4v��)Դ���󭨀���-*��r���U��y�2�Wӹ�<_T�!�k��Ȃ�GU�X*��g}=ǝ
��u Τt���!zh��ٱ���hO���s���� � %�Q�Y����M����0)*,���!������9�C���Y���#�/Uf`�,%q���K��
_� p�=1	�%f�������o��A��[FG����.喨5ɹ�ux*/�->^�y&���誫�*�0| ��NO�'�I��}21��.t�/L��7�k�s�i}r�l;�_�
t�.>%�'68��6T �&ŃW=��I�6`� :� ��s@��x�W��K�l7^��9���N����3�p��9�⎃!d�,��Y��&�	hH���ǭ����&g1A�k��p<Xz�ۦ�����f�=6��|A�A��L��G����L���㛙����ш/V���ˣ:��D��q��G��G ��lr�`p��{�8bs��佯"��x#ɒ<v���|N빭ۖy�2DF�,�j��V�J��v��C@�ǚ;�5u��)Sѹ<)0̈́lk�9=��+��o
�E�I�A�"�3]�5�5���o��� ��yv���{�4�Y.������FIw�
]����[ ��P9 �pⶾv1+�_����èfֳY����ȹ9�E��4����?��Web{�(΂>��FC��rw[I{	�t��>�!���:I��+�pl��)�Z
qy$y
gm��|�����7'�{�ܫ�=؍yk��^��4Ak�YF�Ļ?�(D�6IfI��n&=���!���M�R�p�_��N�
���h����L���	�wNŉ@�qnbE=a�U�I)}�q	�?D���2��L��:oo��?�#vZI�BQ��A>Ƣ����g�$�����Y����\(����h=�:��iq�;�_-��LM���:�$y���2P��l_T�f�y`jy��.Y�S(�*�߳�u2��JEp��y�[\6:KC	D e�e�%���Jlu��1�;�`�K��;�U^P���%1�.�ՋB���1���D�,��O��N��p}|^9��""[�Z
�N�)7��j3w�#$�kf�8�9�bٙ���cVt�o�uv�'�e����hf����#�Ȕt����M�{�3A�vM�a���Y(X���3���%���>�}�����^��rzu/ac�K䥴�����2:D�\j*Y���7�@e���+xQ�+�K��L3R*��p��c5�l??Pl��yȂ�7&����gm�ذ�L�)�I�^-��ʊ�;�F�c�b��ą����bqC���N��%w�;bSo�΢�2�� _�#�d��}GM��v��,�=��ƣ?ë�T���+l��t���?���oW�
� X��¢����+��u��
$T,��z>oTl�)��C����0��J#�O
�vs�t����A~��j�S�:D<�9`��P���wAiE?q��m�I���'0�:Nh������Rb����p3Y���'�N�`H�I�."z��F.´��U��yl�'���������BD��nqS�\&�K�P�m 1��⼊���[! x�X\n���<t^�x���9��pY���~ͼz6RLOW�V4+Ѥ���=��M��N�e�!aUR7xߺ\� ��?N6̔3H��R�%��(�Q�F�%k��I��p���؈;	U�'^����.5���O�pW¯FdN��SXVoϫU>R��.�7��j�|���Wθ���JZ033�$]�k#[�k-��G	k�O�B�XԻM�esrz�|��fB��GPcq@NX��]W���>��|�u�:�����+��|���X+��)3�nSU��d32{���O�e⃘+?�Z�������>7Bp�����~;�HSܢ�_�D�(�7[v/W<λ�R���n�m��M���E]�9�T������I6��v����B�eː�׶F[㟛~��*̥�6O)|fY�A�[�,r�G�#S''�����~j�j���c���"��s��H�@���wk<4� @�~���n5������%G��,�NMx��sW ���f��d{zg�%cI������X�yL��<.t$�Y]��������by��WV�\�k��w{������Y$��~g�2ſ&=��{�-㌰�ݡH���:�͒�I�`H|�v�@��8wE=yTJ$&D����-�D*l�vca5�	��vtDf��e���Z�)��ƚ�'��\������Q�"S>�<K��s�aby��2�T}�Sv@�J%�VC�xn\��jZ�
�6n�8��˥��v�"U%�踚K��M�ѻ�3l/ķ��4ACg.Nb����2�ʨ%�%f�s�ű�w�WR~��`�ћ�c֜�p��M�޾��G�ӊ}9]�x�T%;�w��0j~���ϗ$	��N�N��1a�;��߽����S���@c���.֪7������CCM{p�/���� �9�)�E�y2��5֠Eߠ7<b����?Q꺉�F���v�[��w�o��gf,�XY�M�5��p�x����uN^��D֯E�X]U4�?�����zEv,t��P�������ة�y�&���b��^�����4��9�pi���<Ó���IPx|5o�،9��l��b�ϾI�ӧ"�II�O
���z;]0��0�7ED�'��q�ڵ�")ZSy�%�ϣ�u|㨁!��e*G����љ�4|�G&"j��,&�M'����m�|��8<@��k�0�ܮ�x؇ �s
�aUF"S:�kj�?�� �]�\�j�S)-�@i�4X)&�5��7���N�z��Iʵ�����M�i��):O�{�G���J�A�Ȅ{r����;[�9�ku����6��R�4��=d��:E�ip|�1��{Kfʬ�[�
���.�p�0M��6%��WY��蝏�|&��
w�_��P?��UA�+�����i��Ԯ�kyjI�����GH3s�o�����4Y��/W���:��+M�,W��\-��]�,�ʎdG��3mR�Aq���^����gQ��B0����rڂ�������T]�INV��T�X��K�v
��8�g��W�S)�����}�s�3�����e/�[!ʬM��NE�t�+�������%V
�r{����)� ܤҺI���V�=�?<���ƞ��¥ߧ�
�H�#�{�8W����%~\f>_��a�/�k���Q����0W6��=�\�\��((�c�w���"���GJ�)*~��|Ҙ��cg��~?����7B�	op@f�l�~�S�MUoü�ORp��1J}����z��,N1ٌ7�k�5�l�k��oB��5�s�Ê^�d�d��|�7��B�GU9�"�C"C��C�ީ�QX�c��Pv��+��U�H���p�+8Ƨ����XO��/�	����=G�:M��2��5�o����կѝ���_���U"G�<���f�4�'��Y14�֟B�"�5Ŝ����hO]oڜ3��`�]Cݒ!����42�{[�,���U�s�i�kjq3h�4�{�V)��_"57x�������D��,�3����X��+�HC���?�������]�17���n@M�����u��3K%r���?U�A�8ӌ@_���6Ѱ?�Orq�� �f�3���������p�� խ�N�bȌ�$��KG��~���dR�9��``d,G=#�����s8nñ1E!&�c�[�����")M ������yjU'!�'E͇��>�OM�מ�Oe9S���)5t�:0�>�'J�s~��B(�x ~�AǢ��L��K��cS�/��W���,��H�#3i�|��\bfc�Hz�=F}��Q-g�Ш�v����5s/�^��_�*Q��FIg[��ۅkOˇ���}�$�r&ɊD6m��'�/Kd󆁍�9H��z���W\N�@����q�QM0�"��}�۞��p�"���a�D���̊���<�E�o��IS#2A���W�@g��ӓo�+7c���^�V��>_pSg
AIzd����n��E1#���ʗ`��{O�g��C����1o��an
d���WN�<��Kc4���I|�H�U*����#�y�eX{ID| |#�'�GJ܈YT�k������s���,)V�RW)n�ħ�vT8#,�d|�+�5:7��*Z�m� ��-+�BK��[�.���u�[�3Z!w���)I��]Qd_->ę�뫳�`g�0tRL
a�n����$,��*��_��LY�����Ks��D�1���f�F_}���R��9l�l��^�8G߅4,�6�Ջ�Q�����R�A�6�fZH嵓�
�p�#(�L��Ԋ%�fd68�l4SI�(}_Q�tF=sl�ND���j'��3�-�}�.�=�kHH7_�	g��Rk�C�Yٴ{bO`���ǀd_|i�]�?��e!w���n$nE�;HK}��d1xa���NVXt��cg������\��}.?�Hϡ��\��b#=�W ���@�lI�K�u0���/�	�hPx��~��]}Μ2XSm��A�d���t�h����DNf�"�"q�ɚ��[�v��TV�k�`�\%�8���{� �o��L�Wh=�5R��e��Kԟ ��n�,��X����W	�M��%f��fS��{(�s&�����;�M�1*�e@�7h��� Y�G��!�(�j�"tl��.b�'*�a������Do�Z��=C�R�>Q����#�:��"C�>��7$�@�^�s�	m��u]��G4�9����N�hB&�6؄�"�I�z���5��K�5� ����0<ã�}ŌaTN���:8Q{;����C��n�f��$�;x��P9�iK�*�l����wk�oxB=aʩ���}t��e��2oA:`QZ�]�܋҂!�XG/��)m
nHf���cf��w� ~_ظ�(D�0)��{��uʳ�Sg���|���P)�+É�qx4۶��*�����R7��z����F�XT[!|pZ��I�
�;_��'�]����İ#0Fb�p��E����s�D/t:�ȟt�7R��Y�Q������r\�(��_p����uo1��=q@�-��K^԰���*q0[�
�m�vD8���NvbwlR?cp*�U	�D�#O�E3D� ��_:'��{�/�ڐ'%��-	+�M$leY��\�i�z��Gl���6y��˷�*om���W�C��8E�b���8izk=�?�����g��b�8c��|�+J�D�4��88��w����hXQ�S�B���!깠���2[Y����r�����I��Jы��+����[�)c�/��fP��R��Ⱦ��Mx/=�<2��̡mY����`Y`ICpo��[���>X6x�.1E�M{%��L�����g��&*�$$#֣��-���2�'���%0�Y��[t���gi\Z�_9��P�N�6p�������`��%�WH��kyLŋ��B�x�"^�h"6sf�=�
�pV?�(Ih�A"9�?t(S�q�{j��n�줉d�F�����z)��h`��ҘGAo؜�!�+$��*&�n�?�HXfEW��JB��2�}���=����N�Au�W
궁��p1�W�}|��u��͜�޽h�hD$��D��C�%j�bYh�G�w���Q�P~�#�;(*�e8c�oҼ��W��?�Nn�rF���y��%+���?�]�zX��6�{��e�[%���DK��h ��ݑ����yA�1�N��؆8Y�=�t�o �m|�3`�4]�}�~G��
�k���i�37�'����=�*HR�,P���ꡉ��2JF����ԟ٥i�O'�J:[�֭TPYQ2੄�̕��F=�2�������W�O��a�>�m�.���X"c�/���ocJ�߽ ��䄚�/%��� bYP�V
8.�qu�e~V�ֈX���"E�b�)�g��s>M��N�Q �i�0E�>�7䁿'���#��-�I`�%��x�E��;��}�5L �����h���IyhY4���a�V�:�iZ�"Nywܾ��;��+�%la[��}Y�,g��,bԸ?���5��N	tƢ�����8a�r��	�8A���)�Ã����I܁���2ݭz�؇����"�
�=�>�ɭFP.�恘��(��;�;{{�o�*�dvzq�D����X��
f+G �����T1�AII���A��KD�W*]�a1��#�oU�&8�]����6�P�2�V��J��\� �\�a����a\�����?<����|��|߷������Q;[�a���O��gŢ�Ί8�'��b���v810wA����y���j����b��k�� �$��ʲ�s�s���2/���y����Q�/JrIN'v��Sl׻~O%7�_��+"�i�@e��`^j���=N�w@��=���ta��7Sy!�{�RY���^Kc<��ma�::�v��գ>R���G�x���^NFV�L����֘.]g������P�?�!��aou0D2b�e �ا2A����['��O����0�H�ׄ�ůf�΂�i=�E^��fx"�P^X�
�z������#L��A,�ܴ�;�9���F�y�����'?�!�ⴃ�0TE�K�l�^;�*�K`vl��� �����*�k�����?7�y�D�H%��3��vL�-m�='�d��V���������%lʯ	���:vb!��xú ��\Q�^P�}IH�'�Z�VS�@e��+��xh��w���Y������@��|l4]O�"�l�}��ڵ_����4˃r�x����j:�)n6p��XV
�'��4SE�8�K���p�nO3���q�ƺL�C2sb�eh�qI:�r�ϺH�{0	�g���Ư��&������#�>�S�,0��&��#D�-�\�l��ʫ2��Ր�{�6���d#E��[�=;��w����Fɩ���ę��DF�@��W}Ť�]l/�2Gm���ҷBܻMS�������;�'s�V�{p8�1GP�h]S^a�ɯ Bt7���b��Q{�T���3l*]
<�cn�⩵��i�< �X��f�R/+	��^1�k!�̠���8[(�C~")��������te�˻f�KsC����;ZS׍��/N�����E�-Z�l�{k ������?��b�d���ɏ�Gu���`]-X�N3��k��B�߹�Ydױa���.�nC�m�n��^���Vl�!&�=�Q/Žh,F�!�H��;NĹ�ض��7�Y�,ƘJS S,���NJ���2ӑ�lpGWK�Sd	����.���q�f�T�`��1	����ayo��n�q�ޏr_zY�E����ɔAC�Q^�ryn�l}o�5���S����0�N��c� Wp�v�$�Q}�Z��=� K�k>E�������A��(��>�Yo�܈���B���6`i����#�8S�S-�+Ic�kf��U@�_?x�<A�߆�-LE�y}��ĉ��G<�[��E
��s<hP��uE���k��q�k[�{O�F�U�1<��|1X�M��fS���2I6P�V����*����e��}sajK��]�$U'H�o�6��qNOǑN!�
�Gp�P\��:�T0�Z1=c�h�jU�vN�^ƐԪvi�a:����M/�$�m���dfR��鞒<D����tғ��bw�VФ��C�$��1VYm�WT�����]l�Bp(Gٵ:�e/���ז4/�Q��z�c����1$���;n)��x���Ip�.���V���,7�$/
At�b3	� ̇!	��ǧj�Pʮ3�?�j�jn:z�O�~���a 1�EpgrO���SY��Q� ��E���Cu�(޿<g,��N���t�#ʔ�#�g�ǣE�ߣ���v�P��g@�E���/�ߩ����T�a\�a�-���,ibMej[^}L޻����T��})Y����y�=�]�.�������x�|�|���`՜��$zl�.�=�i�K��#]�&Ey ���7��H[�x�v���77x2ŏ$U�6��?S���,��[qR�H�����&\ٻv�A^_n��ӠHCd@m�V�W]���P�%��G�(���$	Q��+MV��/Y���J=��i
Y�]�8hL�C6n���/O���'�s�A�p���&t6�$W�?����f�n��VE��Ũp��A&D�a?�IW��s���=ʾ���[��GX�'����7�!=��� ���:�n���ζ�l�{����M�UyA��"yh�Dp��<���e[�\N�wL�q.�~?J� v܇�j��xq:��m�U/��w6�����!��v8uR̥����T|�lg�[�>�2v�Jq���i����!Pe
�2}�BӖ�*x�/�3�k���w\��3����8��G�'v�E׼(�@q�|���lGW~��y���$g��s�tm�2�$�
(4b/��L����*
��q\֜/c���+��˸,��q�E2o��.)�-��&�.�C�G��3����5�$Mň3��޺��X��w����!p��S�>nª Ц]�j(�bh5D^r/� �o7��q&%��Ξ�@ _���\=� URB��|'���}�C���@$��1n�����L�'���"�K'���]MMM�Y�2�.bP��.�5��'v��M��d�ɶ[��f��k]3��H^�#��*�x��BF�6��u@��U{>�<����5Վ�!q����Tu�ע%~I� ��Ms�%����m����d�8�A�	�e����C�{+��,	ĭ�Zs�Ƀ5y'��7>}N�0����$���X�MX(7`6��G�,�MId���g�v0��o��Tݩ�C�^�x��R.�6@ֳCp��=`|�k<ó�����qBN�9��;{c*�,U$ufoq�O|�e�r|�7��@2���9��1 ��C���Z���!H�,���٠"T�ˉ��]��'���ߏN|D�:R�SAp���l�Fǃ#����8B��+��U��N[�r�9MN+FI�F���j6n��Λ�۬���|�A��LIQV_U[�� ��K���p��J�u� �����VK�Bg���e��u�	�D%��@*Q>��K}O�$�mq�,k�6�)\"ib 8B�!#�4�e��;o�P4H��{E:�ؖ�N�;�TZ_�$�� ��@����,�m�3�Ƃ�&��7L�?(�荔6 w>sK��T*wA=���&�#O�͖��}�w�v��ۼ�B��T�7K%�LsK���~�)v�F� 1?�7#i�������66�8����b�'�������{*4C�l!6�ls��V�#,i� �~�dP�m�1N�B���|�|�=���ɹ������yw�N�ƲW�s�,#��|k,�U��D��(!�A��9�rl?ƃФ)`���[ͯ�"م�;r;g^Y!�8���t-��8��f�C�RȆ`�$��eP.�T#���Y�.�ĦVצu�����*u+�:�uiӔ�t6���R;.���y)�*G��1ԝ��Y-���r��>�#w���e�s��9����'��X�ݯ-W�> 9ӄ��گDi�½���0cHY���%1Y��\%u%V7����߳�S
��^�~/a5��
==��U�v��!Q�? �b�k����7�?7� ��
��Р�/(�~����s��Xs�[-�ԉ��4�J7�j�{�h�(�QY!��^X�M�a Z&3�bt�+0�F��u��}1��
�DfQ�Kq�ׂ<N0>�ȇ2��k]ᮉOL
�@��Z&�Z}O{��ts��a&X٫�p�r�������
��#�"3�q�4볥Bl%����؃!*Ju2��m.P8��_LR�C���z��
����Cz�[��$؞@��Iw����3Þ$ K��D����P�/�|�e�eg:_����J{�7	{ ���2!�f�Xo7�놥��s 0�D�WX"�-�<��i��R6Ka� �� oO���� ��p|n�Iw3e	D�t3��V񓮆�Nֈ��}
`/P�$<�Z6���|vg���~�Қ�l��nWCU�j���O�z��vT.fP�'>�[h�Ւ��_�wtV������!ÿI���ԣRC�b�h�R�;K�?��a���Ί��и�b����:z��D�Q�R���"����]0��V����(�����!h�| ,����KjXo���:���X�.4��)�[;1J�7,ޑ�Q���y2>����ج���Sy~H.5��H��	P�ŝ�1K�4"`�W��ܞ$�) 䉻lm��9��Us���H
v>5���?���s�ʆ�'�w!���F�+��n|�E$���� ��bp�U�@8}Tj��}��Cy�م/ ����K}�d]2�Q!E>j@T C$g��Ec����.��>$�~�X�W,�v�� F�*������]9N�)�܉�����߄���s���P���D2��5�,��G�e���3�Q�i�*�8���X���s�,6en�ZP�ӂ�i�$�/pދ�$�Y�C?����E��rq���|���z����w�#�4գ0ێ��b@�|�K��e"U�_�V�W���5�qY���KS�Q�W�a5���5d-ag6��u����=��q�z�,�\#s��P�H��wi����_�3���ۊg�����]�뉯����ׇ(�=�F�����h
	T��{�7~v�#�V�_7�PLobD���K���e�j�+8����A��Kc����2��t��<<���L�"�c�C�Rj����F�ણ�����p%25�$��˻#뗠�ی'��wzi
y�sa��E���0V��n׉�E2>���pƵ�~�F��ޅX.���k���b��yƤ-�����vn�Ƣq�͆�����k�9��tI��mu��%��G��,@2�R�#�]� 2h%���J�O�I� t��fKmb��R|�%���|�Dﱀ��ό��_�o��s¬;��/��L�w-a�=�?
�!����	r�$}�V>wJR>bd�)�:>�c .�V�p%���K(�E�mũy�� >�s�A�z�l��1�G
!�a�N�Kf�~��qP�L~#�;{W'�P>}�7>�]���9I� Ig8���c�u�E�b)�l����68��ȟF��u�нNZT�;��S��J����r�1�A�6�i@�����`L|�sPSA]�靱���pY˳�B��e^�'�q�<w����yP��;�c6Ԋ�C��-����v���9�JW�1�\���h��)�L-��S �wc,m��=R8q��4*Z�O��nE�2y���|1=�Dh�]Ԇ�IE�~J�5���w�)=��t���t�����f�c���;w������mlO�?���cѼ�:mK/�K���'�Fm�_�e8]��u���!fs��N�" ��}����NgD��q��M)��^vM0�W�eQYFC�C�:S]���(IH<V�e��`�%���S�$���!9� EB��ݹ�Zɟ��ꕃ{��͟sZ�y�'N��=p���wr/4?�# e���f��S�f��~�����#z@��z�q��J��:6h�a\G:Bm�|����x^�K��zb���?����2�K��4P4뮑��d6 >�����i5���A�h�s�YI��B�ɂZ�Ɗ�h~5�,�
T���kx>=��˅Ϊ"��9ݥM�i�>��V�l�6�	��̰��+�[�*n�2К�����3E��`3a@�9Ų���Њ�X�h��E�I���|���g�U�C��r��B�ϻ�dg� ߅�!��l�g��#2�ǜ1b�{M#��Ñsbgw�"�=1��	��-m��$�n_���M]����*�����o�s�ӊ�`ă#�p�[�9��e<?����)f�U@.(��vք��n�,3�#x���Sm1-Iɖ<�2Ko�,�P������t��s��l=J�/��1Qsy�`Ԡ4����"9�Ycu\zߖi�e|��<�"%Z��X�#%����l��-wg@�n֬�jy_� =s����+.�$�3�0f^�(82-�+����w�]\]7�q/&k��H��G��Aa�XU45C�2#:�`��߸O۞u�U�����Lc�(�Yڍ�|HF�-���r0�q %�` $Jެ�����.M���m�P��;m���^�'��t���Ӂ9�Q~�)%֨4ŷc����(`D��3�l{Wח�6�SE-m-�����(k��P�[Vw�М�����hEAǶ9l�=��h��`@��9��Gm���dp7�HBG�#�a�b�t
9Z �ƫ"����D\��_^�F��QG�51���j�V��w�ڼ��G:��$wȤ�Ƥ$��ў3�J5�?�x�˻���,�¸�?G�t����DiR*k�����(�ήb�eћ��kDM�Ԭ�\3��OO��'��1q�� UY��x���k��t��;?�)O�����Io]���k�B�NLV��۰���g�<����Y�
�|p�,��)?�/��^�[~�;��c��WW8��oyu�p�ދ�<4#GN%�A^4՟H��
�@�D�(�*S(˜�UK`\i�����p=s��]�%����I~)&@R�P9E~����x���$*��p���,k�9��o�?�W��t���W�ץ*&9l?\@�R��nYW^��r���J
��Q�6фt_8��_���CECk<l+��� x���e�e�D��;��A@i��ſP%�rzܮ���->2,.����i%�� vɶF��N?87����X�
 �lKٖ������ �E�!��V0�?��蹃<%̻�"���iL[�}�Ѱ�=]���1�Y�8]���7+-YQ�I�MSC��!��2,:Y�v�Ց�|�
*��J��e~q�ni�ʷ	&d:Nܸ��	���8*Z�B���W��(Om)�E�[h5�)�1��>jK0�(���Cb���}���+�^LȔ�C&�w�8P����\D.6a��\���[����w'.r���gr�ATv1 �ֻ��J���,�m��-��n�� ��@R(_њp�V`��,�a4'�����ڴ
�+֌����Ļ.�\�A����{�o?G��S���ȑ��"�4�����#[7U�~:?ƇQ�����)�n��|�!z|j�J�C�tv��c��$�����FT+Kn�*ۚ�q��a[�F�B\D��!|�T�e}C�ȖhKIle�eW����RC��؞�@@�	+�i&4�ߙ���,��v�(k@�t�6�xX+}���\��Pv���D�$C5��� �\��=k]f�,�!���)�.K+J�&���Y�y�#.�%�RIxF����Y�(uS�q+_M���	z����4~#b}�S����%���wiR���7} ����U9HI9"��пx��wy�\�����7�:��r^eC�n6d��ō���^=���i�Bg@_�=�D�^!�jF�lǹ�]0�+����b_p��-���7^��~+��~\�)&��}���{FW:�+b��L���E�pvly��!���|Ș)�Q��Єq{������o�&�62�g	���ًI���1��j�}yC@�����@�W�� D��|.���i��m�A�e�?lxE(�io��OǻB^�����^�����;�lB�!��`��zm�"b�\��ND׬A|?��x����kt�W�^�l����|ʢZ�s�4�ZjN]�-UT�&�+v��AJ�׀O6�~C�s�#�FGP���D�yK�<w�^��Â�� m�%�����=���P��d��w�yH�ʖ�u�c��U�Ǡ���H!^��I��aI.<�_��:9@$����4I?%[ZļC�G��zV�?Ѫ�r�-@���� m����Hǵ­$�J��SO�w:��?G�B��?kΛ\L��� �F������PA�#ת�\e�m���?ţt�_��9�L7����\QO�8�H��� ��Y��	u��{Ա��6K��`H�Df�2�+�(�Oۭ����ݫ.�R�	gSa;��K�����U��^.5�9����!Gt���3:V3�������7U�̂�h0"��8lf
P����|������`i:cY%�b��t�r52�f�����?ց�1gY%������
>�al�oΣc����To�m
��\�ͳ.�k:ja��2K詸(	h�+��Ȏ��ܻ��x��� �l�� ��L�������O��	s�r�lT	E�/ܵ���a��O�-P@��)OW�"��/�
��-�x���g����3y	�]ֱϵ
{�_�5z��FTO�)����(���{~S�AVӎl�s��k(B7�������C�,Hi��}��D�KԳ�#d�J���f�����g�(6ˉ�?���N�s�g#��'�ڸ _����񋺿}	�ZA�|�wG�ov����Pbm�����2�YƂg�I�l��/����!λ��U({�SK>����!�#�ޖ�4�E<�G$��ذ�F̧&�����..4�(B%�� �@F�3�1&O&�G�����o2�s\ ����\-���yT��j�`:x��!���b�@@�GNUODlp9x!A�l�Y}@� :g�;�RRk	F-�E|���_��'��E+�=�6��۬�I�Bz��df��ЀR&���Tz���&����ux��@���,���GY{cI
Y��б92�^GI�b%W���u�3��ap<�B��p^�p�.��� �Cҿ����1�>��� }�}����Q36��J��&�o��睮�'=f��@�u`�@���q�f��Z�^~'W	������3U�1����t�@�������2�Ys�a��6�tq.�����)6cM)�|�5@�KT��Az�a��Cp�W�pסh` `g�GE����m���2��1}=*�o���|�b���F����0�I��+�����r2#�!گa�W��i-�Uh*�0�!ؙN������?�,Re2Ź\�2��ב��� ��(~�^�V>6�ȕ��t�c� �:�/R.}Kag�o�k{ڃ���u��xqxY���z5(y
�n����Sv-��^\���Q|ꛠ�K� s�v���t��r��2�]���g����:B��{�R	(ko�[��Q��4�����	��x�uׄ�٨�U�4��ss�� ��CAz-O�ѝ�(m&U��)>�zֆ� C�S��# �?G��Bk%�y>���u����C�:�@+6�vf�KE��i�購A~h��2Ym����7�ާ��J�
���>�|�\�4828�WC��u���x�~��ϝ�ʒ�r!���J��fF_7�dW+�i���)����3�=ф��g��L�?��%#j�<��ό�@���׻�F��&���Y'��-���m��^�d[�;v��}ù6�Zfvw�����M��Ǖ����(�w�lbқ|A~�����IJӕ�40'm���.�sO��w�C�ë	#�7�񥁭��~�cc��|��y- MkC+�D|c�Rd���. i�=:��?ݜjs ��̳h
bu�� ��#�1gF��HoҹZ�8��2X�@�4����-���Xw���!�P
�,_b
����.p>��G��{�3��IaN81%ë*�v[.cX���32u��8ۣl:Ć�����uo�0�R�Z�5!�dX��7���x�������|I�0Y+� #�)�7�l+��6���E�4���o�:����T��c:�j؜>R�º��!,�mK�v��D�,O�=̎��M��Ashr���1��� �t�|0���p59=(O��|Z'��݄" *\��������,�+���Q��%��+#8��;��Ħ��g6Zkac�Y�4�\�{o���OU�5ߚ���g�� ΁U�`5�~m}kc���.A����>�P��ײe�4	����J+��FUg�n��$r }��8�x��}�R+���9 l�G�U����ᠻLB�0��{�ן�vi�-�Bȑ<�O| �h��#?j�ęh�������1j��=!����%(�t��5�}@�!,�gw3�
�2u�	G܍��a�{h>`Y���,D�L�����R�Z�������Y����<,^J�U!j��֒S�s-�8���(����n�՝5QH)9��׈��B�H�)r@ ���ʻ=�		�j� 	ĥ6���ʌ�H��w�Ī����ORU7�ŵ3���1O&���(��4��5��i�6����bꐐjS�X��~d�/8`A]hٲ�u-@��ӡ6�*�'r������(z���������Yk��J~�T�]��2��w��D 	�~'��Rx1���'�t3-�12��JX獩�mz�⍲|+��~��|N{g�3���@���y�2������VLP�zl��&��!<�r�2��:aN�)�ڊ���dBj�͵5�E�Z���$��&�`
'���1�n+����<6��ә�������j�ʘ&Ք��V��(C����K�@��ѫ9�ꂩ4GB��6_��F���ѡO$�*�ԽOc��A�f�$�UF��T������;�=z=�<2�����gÄI �6�Rɭ��1����	��7?�:����ά�!xn%5hg�	0P�d�q�X>0]�6�ciQ�9C(��"�+*�̵��)����Au���9A8"�^��n90��T��s�W"X\�{��9b~��)�Ԃ��M���r�y���vv�;���U��usnkz��ڑ+��u�G���+��@m���N������.�޳�~1�+)�n�,Ep�Yct�.x�ڏ����	�O��j2L()l/\�H�5bB�/�3��������<����k�5R����C��k�@�=����ڿry���飋�bd���7����{:=g�O&
.L�<�['MD6�'�&���^�uEi��C��i`-����z����ly����"B��AI�p�K���9�qFg�������I��y,2D�@��v�+�p�-bSQg�3��-j���e,|�>�)֏���'7��^�3@S+\�ᥟLB>��C�/�kj�2��#BD?b�b����w�oZ�����&v����|�LlX����𻖶1 Iv�,�c��JK���>mV�1��
LA1v�`��>ݷ�)z+��ϲΫV�S1 ��96�_��:�2EAu���p����)I���#eS�S�lM �W��DO#��se1�A���IǔM7SBش�'�2�L;a�\�7wp��#4TX�P�֩Y�rL=�dQ�Z7����y4�`�n�߲��)�3<8�9>���{�[!7�i!y%O�O
R���i�U��FHi�Ma=�D�x�r����D�|��Ｓ �KYQA��3>Ϯ����cU\򫤄�{A������9����ۺ�.��ŰM c��vf!(��Nj
#�&���y�A���L�1v� W������\�	�t׍Vo4Ww�_�]<�s6*�.t���ù{��<�ק~8N�t����T��o�g% ����5� y���f'��-���>�7`/?��b����"��@
���4A���� �|t�������k:\�!�<Q��O	$���S1��?��E��&�Bg��ֆf�u�#����B�oiP� �Q{,�����Z����z��	�X�	~3.�-�'*��2+��V:|�zc6�4E��N��_~�ot_��x�i�1F�����e��TQ�}(�W$ \�����9{A��C�-�+�w) ��>�%�o�e�I�w�վ�Q�89G��D�#�CG�N���������{�Nm�|"�c��ː��P��|�#��){�I�b̴:<�V&����7�(ۑX4�����C5��7�Qգ���7�z���Y����E��h�) �|?���W�gQʛ�hI�׷m�kJ���dCJ[q�g�7�Ͼ~?N'�~�p��eF<�]r�N��{���9:ӻ�q&��מT��A@��kz@ <��0�9�|8e2�M���� �U�XP��AƂ#������r���3�'n��ސ�Ғ-�s�!��핝�Ar0<����-���(N�.w`����[	��h��~wm����pU�MU_A"��Jg�y��?��c�з󗐝��u�Z:z)D�7�@q�צ��M�x^olkbH���B-��`~vY.�W���&�=*RQ�b��"�����4mB�b�����%§�<������R�c(��Iq��l�c�5P�صV1���x$#����%������Y2��ې|�Tib
7�F��H���Q)a����S�W��`n����ƈPa�"�%����[c\Y ��\"�V�,@%c/&����Q�jI�/�v���<_I�Fn	!5���ODZ;��F)�ȳ���伆U����a;��|Y����Ư �������D[�ٚD!؄�#�
�vկ�	lLD��7{aJw�k��l��'��S��O?����Gg ����HJ��N�������d�#z��Զ�R��N�8
"���U�nJՕ�2��Ƕ[z<��xY�f�8s|��=�o+k} �F�bi:~�#"���˵���\]l��h�[�4%vL�[��¢R�����{�9��ӥ����=W�&�;CzQf;���I@��
��h�H<@���È#+���R9�h���!`�T��ehp5T�o�L��V'�L�o+��5�D�<������4zb�T��\((�WPA�{:b@cшS�`�{���V Y�-Wn$�;LlV95���T��������h5��@V�F�� Tt��[,�Ҷ��B��v�-�8�J�ʜ����"�c���E��+�H�-���#u 1�FM�H��˂Vt=��9�z�'Au��8�Se��C�ƂKs�3�����̜��łjL�'�a�`�Ǧq\�¹r�Ƭnh�P�,�x��>4��<U�'�᤼��?���w���؂��Ǐ<���7�6��K3T���\�V~Ź�	��6x���u�h��P�Q@�2VJO�:UC�kJQ�����K#��5�#��/�8�c�>�Y�?C�&>��_�΢c
0P�%:��#�q`�D%�U� ~���˸�q����a� �g�{?��+��5���-�1�)i5+��	 1��u��Cq�c����y"� /��eXã�ˌҮ[O��)��V���su��x,OVw�E��nB�z�]��Y���d���2���Kf�	y�0%W�S��}�㛬͐���}�-Z,%L.�v0���x���ͦ���G$6���jL&7���l�;P�<Q���9z����c���p�g�\X92f{��U>GϮlz1P����ߗ�Kx�<���K��4�߾���NBc�u������KAX7r��c��!�ٶ�^����X�F�t���l!�4�k�{���!l���GBwOբ�7>"/���ő,\����ԙ���8q�(��ɴ��Wk$%���H{$�*1V
&k_��"�m�z]�;3
�`m�<c!�bA��˺3j�f��!J��(sq���wj�T(z�uЙ}G�"�X(X��1ǉ�#�$}��g���\2�XJ��Ot��;�T/�����6�u�Y�U8_g�t�o���_�2>M�c��]�+L�֐��}K����7��s�� ��C��ő˪����*�m1��wy۩՟�s]�Y�Y⬎+OR,�	�L_� �� ҋ�Ͷ6�颷�<�Ur��4�bŷ�k�3Tzm j���g�k�T��Fh ��Y:Q���������K�F��ߣ�z<��b
��?�o0)�'���	1h�S-~��֩]=�*��#��3x��|jr�g����WM�u:�g����AV�zL<�\�,sY��g��Jv�%���kz3�JJ
�'R�?�-Ei�{���(N��^�C����W�P/-K�:�{xT,�^�����h�,�$��4���+/��-+��<�3u����ܐ��\UOJT�e�Δ�DU�\)��!�j�0�(l�:��X��F��p�*�����22-x�'N�"���A�F|*QЈ⡈re&QJ�V���c��z���˽�e��o�	0�g�&W��2)�q<�Z�WL��ܱ����	��H���Z�p�u��_�B(�\/��@�`�D�ZG��qz�o�۟�9��?p��̛v��hpH���b-���|�؅|�C D=v���q'S�Z�@q�<_�=B��Z���_:��>���",J�~Aa8�i���~9�!��'g��P}�V!�dl�����J���}�Q��lO5��[�lҭ���|�5'	�ʯ3ۀ�ɥ��t�o��\�z� qA>�S�(r���{�o�߾M��`��0��E��3�@�Ee)ʇ��@e���(������N��Rf����i�.1��D�
p��`ޑjx�`�=(lZ׷�V��c^8M���w(;]�Բ���S��[�6cju�j��F��j��� ��K�,���ؿ=Q.O�[��Pv2I������t��n�#��ƨ#|��G��\8b�ּ��TW��|r�7X�)���~������@z�`�wiM���}%��=J\*�b"�L|UX�t/�Y�B���=U]�%T�*�NQAN4�@�1��ڿTJ�D,�o�z�twl+[������f�b���דDA!���f[=�~��(M��+R�A C?�;FnS�j�V�i�q1�/�T�.�л$f�θ�Oq���Ӵ���8�Yx�l*!���F�A%�0�qtD��(����qAi�b�q�d�*ݗw����N�e�<�*�
�y]�chU��7l�~���03�6Wqf��Kr���qL?�_��VR��T��{�U��֤B1�)K�UT��N_�8X��nwU�E<Q#���p����v�Q�&$���4�{�r�:�U��)�_
��0��W"�Ż�X�%�#�J$X�3�B�7�GS���П��p=�L�*� ޮ�PX^���2�پ�����$3���TO��p ��B|D��8��q�ҋ�V��|���d��������������}�eg_A�H���#���+aj�&j�0��P;�|�������?�(p�iK�����Pc�u�~v�+��Z��n����V%�:Tr��i}X�z�o%�@����ck��x��p�O���Y�'���`�@����� Y�|�����Tjg,�Lb�9��n�^�P�/�"*�� {�E���������5���]�t"He�Fk<�+��OJ���>U�{��͝�`��.��k�;5u��ZCu�RV��[kzH�@�Ё
]��1yTVZk��8�v�Cu�d�L�ۧ��մ�#@{Ǖs0P,��p_��-:p�ΚJ�J���y�J�-d��Kbč��u4�����U���O�q���E��L.���e��
P�1ʎ�X>)�{�Z5�j���7��CoB�_#.����.�NZ��/�<�]��n�@~\�s�ʈ�=~]�.�BO��n#V��7,�,X�be�x�<]V����֯=�-�{�S����cT=#��DYp�u��ca� 粼!K�ڃΙ{[�3Rz_�bx���ǭrh}7BkS��м�$/��M�PVZ���ˠ�#�sfH,F���ߺ�w��
�໖�)�V{p��w�	K� �;�$)$9�i!�V?}m�ݷI��U�B<��M�I�4�"��	+�T�\�d�,�����F�l���F]{��UeEpS8^�$��끈~�Z�(�Mve���J��,Tzg˥�ؕ:�A�w�a�JJ
����a��_���F����ʰB�>,Ôk����
�R���V�|�ɾ8�Y��TXWUv�S@��������{�ab�3��]$������Z?���AG�~�K��]�y*Y�Y�(��n�,��� 哤�Dz�C�;��I���[���M���a�R=e� ll�`J��A &K�v]�)��*Jv��s�-���.3XD;�)~�t�Ď:X��+��i������U��<�����z(��U��Y�uӞ.YV~[��5�X������[{�����c2%t�<�F�<�\���J��I���,
�*���H�G�(e�1c��Or���h-�R�`���>�?sa�L�u�&�Z��iZ�q:/�暁Ӥ���6g�."�gs�������L/�B�8����8t��2w/�ue4׀���X$B�[{�����O���Q��1��q��������2�հ����9R�h��DB�������T'b"�昮-����pa�����^5��#���7d\�`q' 8�Mчf��Eu��F��m�?=��|ЪzO�!�[�L�,�;�Fp�?���ĭ���"hzCl�aD���t�{=�!�DY[mSk�]�t����8����=~<��e���g�;��g�7�RL���.'�"������̅� �<�	���}��#ć@��X[�=�6��1L滓Q�����_ ll�d������q�!�����{��T�3�� 7�cՏ�߄��Z�#Mz��c@ê:G���@lߝ�աJ�~�H'�ǕAp1)�����x���:V?I�c&� ��(6��6��~_�T���w� �WD��M`׏��b�&~��x���2�:a5V�g�{@�~��.<���|��2�f�b��J���O�UƜ�q{�݀�8�̢��%��W����DyU,s�b�������N�ur���^lzw���8&QJ��)j�M���BG�������Ly�m�B��ʵhR��������n�|��N%�(�a������_@>�[�-�]�����Jd��ǰ��u}��L���Ef+u�î7N�L9X~{�塖ګ	��
7��u� Rx�V}g����Jqq�ѫ]�V;RDf��������:�,������\��Z+�o.��`�LKO�:�J2QRά�t�rg���D�X���8�־�.��>���B I�Xy��ԈC�z����~���XWS����e'�0j�	�ZIm�R�����G
�p���=�Cu�(�u��`_=��<�HBy�5I���H��`	�FUJ��$w�#?�|�'*A���EU�P[�F��vjC�0�&���4��u0�u̬�o_��}��B[u�� ��(0��<�VU'�h��$�(j���
ei�W�6�9�&`�%����!�vA�À�i��2�H��7v�6�'?�jlVVt{��v����J�d�+�YS�(t�tO�M\�ϡ��� ʓ�0�$�D��#��(�ۃ�_sN��ǜ!�Q01��==����nshZX���F5b2�<�C�R��X������hNW�� `>X�I��s�+ƣ$��:�0�(!��B[I5RI� V�I`ψ2�Y�G^
����S����z�c�d�)Q���Y8�B��+k����@It0��S�����d�_΋�m��8@?����϶����D@�y���ީ�2c(�����}�����ܙ:�q05����?;�]x�u�����i<{˦�.3�m_��A1�./��5��Lʎfn��k$�^}�A�Ğ�&6˥�
gD	ȷ�u�(����p������	D�������bд`��y/=��f�F�P�|gW��5<��q��v��"����A������%0������<�HPg ��d�y+�y��vʢ���-Q�`�f��H�ŀ9�v�eW�u�n�A:�d�F������
6�x�/t��E�z��tY���i+i|)Z��ZPށ%`W�_�3�%����=��2)���~�X�X��t��@�`G�V�u��w�/�}�`Q��`�§��I�b;u�ޛ��k���d��G��w������o�ϛ�}4�Y? ��X�P�Ś��?g��Y�i@���E3�s��?����������v����VRG}�u��S@nv"���@Ӳ2@E��5J5M��k�e��,�3�3}�!���-h��h��"��\���?�;�	(�a�F�BJ&�vL`�ZA�ڎ��� ���2Y��l�����x(�6�p-u��-���'�48p�
�褘��Q���5N XJ�>1Ա�U�=1"���"���Ã�,�<;��떮�m,��,Ga!b����Zjh�T��\g�-n������FKM�ϸ��驍�<��rŘ����FU�][I������������<��|N�� �p�+�;<��F_#{��]�lquGW�
��K/>@�����b#��g�.�+��Uzw�~���%X4ƫU��D�; !��FGdZ"	��J��)�/�8��O2% LVl��,��)7=���x�#�^�(��H�����ϛ�OX��8�
)F7k{��. �=Ir�dٻ����X���JL���ĝ���+֓�Vff*E��a�Ֆj���V?\J· ]��By�T5�S�c�vyTg]��W0/�~i��3��V���ʂ����@�lH�eH�3���N�n뿐/M�f�C�0�;�e�!8=#<.c���nU��t�b/�Q�u���*���R�?�(I�G��D#�Z��-&����s�Y��S߽4��m���N��Sbq���dr8%���ͼ�6':�!�O����}�(R�����{�L9��_���&��MB*�J�?;�m*{�@׊�.���2�]���MX�@��%ނ��n����ݎ�:��`:�hSML�G6��E��.]�W�:L��qi���`��R��� X�-�Κ,�-��WZVz��*b�MIB�8�Wb�;/���q��?e�*�C{��,�>m�&�Pw�z�G�$��.�Z�Li�]ݶ�,a�k+���\�)��T���]�PC=�?�qz4�Kњ�k~/�I��A�Ύ�).;��a��"t��u���L6�t��r59:��c�<�*<-������-��Cg�H�d�=c�ɇbf hP�-���u�P��Y��u������4��������r����$g4�QO�/b?"}�hlk<)�)����:1��U��)ܕ�;*�L��ϐ�;������������*m}�=>-�L�Y�����h�����aO�`ۜ�H�}�@���;D]�b�TÕ�T6�9{�n)����#@f@����3���gte�|:̸~�H2@��\��;���!��?ʎ���\�����+�J/�"*j�U�C[R����et���2�u@��Ѧ�CI���V�CDU3`�.�0��+TyI��_"c0�-����<)�-X���z���� }���k�o��3	����]�\��̜����5�@�p��5�*;�N`�f�Z�smX�ø|U�I#�7��R�w���R6YU��$�����+�8%&/�<�C���cDt��댁8&r��'^���}
4��6)�!�j �s�:N��O|WFCFy�&�}��kBus�&������ᚆ17�4_WO5��Ft�욵պ�?���i<2�L�
l�*ɻ�����'=n8U>��]݄q���c&f]�vʝh�i�[��3��|��	���{���k�9*��N����at�����?
�hU9�iuSIx��b]��{QMa90���ܑE+O�	6Z���>yI��A��nZ�� `�4���{@4�g�gM������G���Ao��<v&ؐ��w��IO���?	�L���ٞ��ř���>���䥔���!d�ю�Zǌ2�>��G�W؎�̵��-��A�R}��$�{�Kg�%��b؆�˲��ٶx 噊��s�(M�:�6�Ώ�XMFi�����=a��E{����pB��Rp��%�#��8S��l�s�X�BΫ����td���% �>[~�C=)�L�`^+be�-�')s������X��i�v�Pui���(�oob���e�iw����	�*�5[Zt���w%�WyPsh{> H}�<�9`�@�]%��r�nyih&'-���?+	�s�1N��mu8�4�&����
���+;�Z`Ɛ�mh�
��O1ns�!����"�~�?7@�w���w3��A5�֪����&�Mz��?�`�!�n̡�#�9�Q-�[c/l�q��l��Vo['��/?xSt��Ǣ=J�)���VNH����W��4����t��yg-}��6�s���0�jNԟM.!߅��oOk?�!5k�%�va_�Y~U�sq���0X�K�;s�a��;�qZ1
@__�#~��52�n�8h��w.|����N���'��5�p�{�aџ�OH�p[�=t�c	�8y,^[%@�ra.Vi-5%--���0�n!�H&�R�7�	Wa��&R�h�t��>ճ�h�O�A������yD���S,�~�@������W�0���Q����S��h��d�ƫ4�㸨R33Z�.�]0c�A5���̞A�֯�� �3O��ewAx��Z��J�Q�gJQG�s�h��d�R����S�{��1�l����Ro���jG��.s%E4_R�qL���A���Y9fC?n�R�݃�'"t۰# �;�ؤ�t�}l��܊0Vh�����į{�oH|��k�Eb�����9Um��$����\�Η�U��Ly��	U#�9C���a��I����[hq`hQ+n����\�l}��8�w@�,2���χ���y�e� �R%���~wШ�YL�2|z��|���x&t�C��WgL�?�d������'�^�~7'�z�@�zf�UO��L��}��:��t���eA#��Z2~��W��a�@��	���E�������7��v>(�V"�B�d-�0Sp��}_q*IR�A~�K_�F>��Ǹ����>�ۧ$�և+��$�h���W�_��m��A�s� �}^��\Z���Q��OH'���,������E��컋-q�����t]��҆"
�+���LN|�UǑ�!+�H���b��n���?����F���z�����*�������Gb�`�c�5�%vϷ��̖=k��ye�%���w�	�M��'��~ն���>���� ������M�
19ȗR[{y^��T<-ѿ�O����NZK�a�O�U�w`�FY��N�D.�x�xA0�$��:v"�K�/ ��PB-���]�=��%�ף�mY�~H�NzS&¿P�[lii�(Q;ߎ��OS]$�!o��h)��whs�0cx�6?f���!6���*��[M���j�X��bJ��8sH�>ZG%l/�R�$2���X������n��bJ�b��������顣�@��Wʍ���9rat�W, �*��N��'�s�+ ?f��>R�k{�Bɳ'������B�bc���`Q��|؜QH펓^�\�|�׳7�d׵6j�Gb��僴ꞞG[xu�[jo���'�00vo׿��cC. �廩L�^�f�pj�yo��φ���{F�zǩ�eg����5_��lq��xm�[M��A�2�yo�D���
��(� �_�xL`��`�ae8 �<�a@A�=P՟z	~�C,dW�P���y]�:⪿vֽ�R��Y��p7D�=1�풾�V���F!��a�	&V>�%��- �SE'��{s� ��O`20:i�	����8�8Qk��Dj������2УO0��g�Б#�m�s~�l(o`����+oqϢ���;H\��vP�"���Ԙ�d��gүy�zI�0�D��o4�A
��(zL� �wg�G
Ⱦ���1k�ƳL5no};�;�����",d=�x�m���h%�~>&6,�"���@]�����'p4����KJ\��>�m�t�C�g}^�@�;����Ff��d�d�$+���,�X�x���1���FqةH4_����GUi�#?gfȊ��a�"�P`��@a�h_�`F�G�%����s*j*�|P����|�=.9��C)��#��ː� 0���>� �N�����ֆߞ��!�6�J���.�oة�;W�Ē�+�'����ѹ�]���ʉ��$�Jm��8��4�o#���F��_�Ǝ�T%W��WLh�@ߚo�
�	»>-��j~t�(���ƖTu&����!,>펻o�ނ<ȇ����d�e��]��iD�ڝ74��X�8F� �1):c��1����l���9Q�Ķ&�g�5�&2�4���{���9�8���c���q�# ��2$���UΚ�A�?��=NZ����Nr��2����8%��9�����k�/��Q�z*	��xo�H�̓��O�и��}�P�Rd� j�V]6)C+z�`2���lA�7M�s$ b��sLw"^�m/��/��" �����v�׀;���Z��<}tUʡӎoF7ߣK�;-�4�N�f���9w�g=�ܤ)�[}�-�,@;Ķ�xX��	M�$8�cp#���]�R&v}BKXv�ћx5�J�v�|�oՆ'/s�ՀB ��RR��aqK]&6i;�t�ʞM��U�^�A��H<|$���-IvB�m�Ⱥ]M�W��#yWV� ��T8c��}�P��*|�h�hj������)����8��ԩ�3)XRe����k|Q<`�<t����,H�L�G��t�n��&QMM���=y� ��F`t���D ������HG�X��L5����
Ŵq��p�<�$�N���CZ���PNa.I��F_?��J2M��ARf��&@q�7Y۸t���%�S}������b�B�R��p��E�xCCt?�@p�s���v�9k��KK�$��Y�Uո󍲄P�3�>A�	�タ��H��(��F��h'a�/u��Oɯ��'�3<_N��RU�OgV�Q:�X�qM8Dur�!��;CM�>	EN)�B5�]:��P���8�63L$bn�c��k�x 3�a��w`��x��T��Z��lh렩1���=V�bpyu�5�V�WIմX�kzdV!Z���iJǌ_C���-����Xe���{�����Nl��L	����oYm�O����	��g�%V��@�3��v� y���]���T����Os�ߨ��F���b���J0�7���Q8D�+�Z>�B�5[i�R<��.��P+�\�*�E)y� �\��s���Լ�u�?̩&�C]aQk��T,QϠ�X�}�ZZK�({���Ma��S�� t&M���K�5�n;#�h�ri��n��*��K �t�-5��Z�(af��?��J��)�,��H�ۇ&$�鈗�O�3����t��f��x>����0xb',H������q��;(�!���\�A��x�l�8�L��'��s�H�eWk���֚	��%h�����Z!�SC�a�Z8kw�}ˡ`���:�-�"�W��-�a��#=�W�-I��+g����.����a�e�;�O�ç�E��I�m�.��?� S�y��6�;���7T�����S��#��z��ecǌl��^ҹc�>o��%���n�
�9D�,��ݳQW�Hex�2��n��A����4�L�(0����{w���ع'1(�ne^#��w�Ш�JA(�.ف�(,�[�߮'��a���� c���x֚�OLǔ>�(���������NE|oPbe�!��ѣ���Rg�yC�L^��F���L��&h�����?"�� ��[�|f�)��o��}*i�s���2��r��?�N�y����C��4����w��J���`NC�m�4s��R����K��H��]�]�J,/�i}+1�ۚ��?x�qB��5g+"���G�D)�iI�o΁�,��>9��w��@>[%����D5毘�����!�ʫ�ݯ��c,fcb^���_�V��U-�iyj�j��1�Z��|�{���-m�(Od��r�"N �q����uiH���x��;S�ᙺ�c�����g�� $�i�Tu ;��P�
WIgK�H������4OR��g�I�2�B�|��������E� ��dy��m�\�x���>���Y���$��y,��v��1t�����|Y�ұc�T�L���m��ܹ���t�쳭Tf�q�_��CYn��0y-�o�U��U��-�2��#d9�穢n���+�-`����"�-�5�2�+fȪ�W��k��v��f�F�79�5��KN1_^��Te.�f��mT���m2�͆2Ծ����7�}8��V{�F#]��;�xکiR`.�]
	�%1/4^������/����'8����n<���'4�jq�y ���,&�����)��hmo���Fpb���h���癓�������?�y��HHz���NF���#ut.�r�\1R�T\��e�yA���s���!��uh�j4µ����I�ޱO��X�gh�e���˾ɜD���+a�E�����ڢr��N�^8^y,\����lMڠ�k@�*�����rD���*<����X'!��5ۘ�:f�Ĥ�'`���cSb����~���]�v�e����ʏѾC�]
A�휌�0R5� ��(y�ѧ>��q���M�#y��l��w��_��_5\�RJ�a��|�(�ӄ��-�:T��hzoF��y5�UG����v+��>,k]��ɍ�`��"� F�P������$�����|�w�V����4���Jjk)M�\�o�<�^�k� K�i�!���/��Hٱ���Y�S����&�!Bm`���U���+���x���>��p���ʪ��T�������kX���	��ֿӤV�_�0|�\�nq��r�㇔/�h9_��	�0��M�
�Z@�è[�J�:J��9�wJxC>�	�Ua�Vn*/N�[(�~�1:(�NS�(�2Y��/A�G0�XR�X��~'>2M���Ā`���p�J%�S㲏�ɝHf�Յ)���o�f��Hph��f��lx�,���.�����צM�:�;q-&���W��nwsQ��e"�e���H�٠q����(e��ַ�wl���J��@C����
�_��b���৘�S�����ךLC]-���߼9��5pLI*��Э���W���k��f݂"��0~nU�98i���	��f�W����"�_���o4�Bt?;L��a���Td	Դ6��Z�f|�L�+p�~eH�R5�9@G�ɱ{�Zf�%I�Lk'5�|"�
G5�����*�i-��L����0��
ܝ��	�G"��	�V�<�[/���Yx���� �LɅ��jj#��/z��b��.�&��o�3��E6�.Z}bsp�f�2�1�r���2ž_�B>I���<}�m0���8f�7p/�T��ӛ��m�d�Z��}N�h�I��͒ר�.jf���{�,���f־�9C~�8aD;����K4�l�e�zhl �xɒ
��~�0-U �W�H�d'�#K���		?۫�i.?<��<�~ץ�<26i�-�� HOl�j��
0��~h������﹖8�oE��\����U�Nv]kb�9�^��	����EZ��A5zV�X�v�*Co;Ud�����m�wB��)�0Khl�+��Z�'��#2m9�U5�F����B�~-��C-��Y��c~*�Hڹ5�/C��=�VM���bOe�������kq
�J�|�$�sGu���lmĪDp�,�}Zm�&�dMe�����m�x���A
�
�)�/h����A]���Ō�i��qH`F�rs�mӳ����W���� 6z����9�_�s�g���+|E���\V�\�}"��K��2�v���m�����y̕���y�a,wu�C̭�>�NY��ч��>(w��hQR��$���\$4Mb�#*����&���̓�YصsV$�Q��,�A�7@N�b�z�Q�堗0p[�|�p�����<u&Y��p�̝E�߸sP��� a�$��=.#�q�C�1]CQ}�1�E�G�����S���>qJ��>o��	�lF�����w��U���;�W����qs�j�
��[]��a�S��Ei$O�w`�������t`��!_'B�e���M�6S��Gp+�^@����yd�\ �R�CF����A����&R|�����l�Z��͓^��b����5�r%��	�P����h���+��OT&I_1S�!�O
s1��g�f:#^�7k��]�QE��+φ/�dp�'N�Br�g痉�?}���X�"�A x��5i�X�&�����������\����;7��w��j��y�0#��	"
%c.N�<#����u���O���4X>V�$Fi;���ԗc��3����R"ֱ��/�z�V6�B�R���F|��R��(��;"�F��c�Lρ#<4�&�(!`m[���e�_On���s��^�žmX��dz[tqK��U���r\�2����;�B�'7nzx�B/��\��P��u1>�i�-�ðM���M��d��:y�HؼPȤ<o�$X��㤥`�����ɦeyr��^#*ڋ~��ȝ��{�{��Pn�#����oGoS �>�����s6�2k*B`�=q�=z3t4����§�t���q�WA\�P�h��� ��0����2߳���/m��x^����k+�U 8�S�5���
��__{�f5��Gk�i��0䂙�"����/)��NJ|���@v���Q�����q#�c��v��?��k_��#� LZ��'�'��}K����-���g�U���B��G��RM�W���߆���� bd�e��9�m��V5IRt�t�w�X�j����:������d���!}��S����YK@��e8z��-�ڀ��?�]?�9&ʁ}��Oz'y>v���%D���!?p�(�w$���\���M�u��/fk��F�����"�8~�/����ұw1g��?���L�Qf��7��HkZ��Z���;]���Mo!�<���U�� ��޵Б�Վ�ө�D"rn#g�έ}y�߰���WE�3��P �$��8{~zQ�O\��]�����3�7�01:2S|�9�r�︟���g�7���?�t�J�:W�\��Fz�x��%���\�_�o����R�*�P�y��X���/O�I#��s����}�3C�����O/{E=el�d�j_��d��� ���M(T�c|��UC~g����@�Y��� �Ƀ�T����<����Lf{��!��k�;�b��r{I�]}0Z�G��1s��ռ�
@0i����:iv�>#9�z<@�9�d 3z"S8K
�p�I��+�2�o����ߓZ��t��چf��y���M���F(~_���1(Q�F60S^ʞ�1b�-�3j,_0`���FB��Qڒ$�%�^���F]%3�[�N�B���ﵨ��&��>���~"�3j��s�t���] ��e$�I~aq�ݗJ�%�?"��z�mOl'�w�n��4r����J)>r���>p���0��QI%�\K*0A�B3����Ǐ�Ͻ�C�p:
�_2\!�m"D��WW>�ra��>GoSl��xr�fHJm�e��W��&P��ǰO������TvC[�p97��?�O;()]��H��9La��Wm� F�ym��a!�Q#��a��_^x�.vI9�3�����E8`3b��Is�C��yy��HZ�{?���<!�<���#�f ;���Kؒ����F�O��=a�g;cM���e<�{B$����k���̲�К}�3���S���E�x'@d�J$<;
�"wx]`��ų����k���3hƘ}�So�oI��P_O@����q,�ç��Y`d���aO�M��"�������ɴ�2�U�3�.Φ��_�x٧��R&(G0*[��,Dz/wX,��L�jq냂�[��V��ciI ,���W��N�~ MX7j=H/K;X��/?�s��&֫j_�NW �aU(�Iĉ��O�ZAN��<��7be\X.����ʜ��ƺ��ϔq��Vx�+hŠؙו�H�\���ƫ��PlO�	F�Lj��(R�Y�׆+-K�w�/i��Ud���U��� 7~�ݟd�O녙��OxF}>�G	�K��0����9�gd?�9��ء��0�&�ua#��L�~�R�J�UL��	�Z��ɹ���w�B�AI_�Ϛ�!^X����zx�Gb��W=��4�G�ŤMp�u"��-��Ir�E�ӱ����O&#��tً�v�y���l��;�]�E�����Rv*��<FMf��{��SӘ���H���U鏽���{�����8M�Y)x��M�H�CZk����./��,�zS'Ux�LCI��
��>v��@Y^F��6��玢� f���š�.��9���Zl�>�A���
�DE���9-���س�m+��ۑV�r���񇅯��+�E�QAUG���>�J���������Ţ����������N7���PX��Ű��ry^�BxZ}�Gu� o�����.�{9�	Pt'��1�q��^s���7�� �S��S��a6c��_ć�Q*�X����P��.�M�QNo)̸�/���V�	��j�<?���hd���;W@�E�5�RU4������2�)$��Q����߅+>�X%h��ױ� �����}���q�S��5��E�[qm�������8�/�	�Ϛ�ƚq��pL��rP��h���Y���(@ɖ��^���ޯ��L�V5�pf�"˛�,�l��-9)�#���B���SK����`�%}���k�[��l��2YH�.e ���f��� ����a!1�H)�����y$Ɯ.�'��&_�Y��������Y����s�����_��-�{�K���Z��nԬ���ю�B�0��'���/Yl ��h�����9���c�K���R:ʝ�o��)�V��w^!"л��R��Nl8]or(V���)�X�)d��$.Q�YЊ����f���%a$SOF��pP�V�&�ϰ��u����ߍ������{"rZ�>1>9bN{�>��q{}{�Dq��78�7Ix��D=���z�Y��}�A)����[������6x��
��w����o��62RB�>Aӏ���ٞ���Q��K{1~Γ�ݏ�W�ةP����E��PcԀ��g@�?ߠ5M��y`V�n���l2Ŗ:�fr�q�<�]bV�����1�.�b39�]����7���hr�.�W��=��?����1�`5�9P]���u��#f\���U����S#�w��(��a��e�|>�ǲ%�T����@t�3R<�k)2�� l牛$e��8;v�u��C="6?N>�4[~;�! F.h/7^;5v~!t0���aW�������,���m ��k �U��9�U�8�,��#�w��_ �j, �<Wz�C7��_���%.q!u;ya@eM��V8?&��@��z�;M����I��Y��S�-��(�-}�*s��L�#�q�cx:^2�v21�[W��g˝&�=th>���q�����1{���P��{���qG�i㐗�,�[VxZň�v�VKf�i���«uM@7�6,�7�C�B�iL:�<��;k7�m
��E=�POq��i�cK�9�X�"|�(15���Z%�����h��wh��r�pIN��^>T^d�z��o{JQ'�%!0 u�<��AR��>�O���.�Af�8�Ng���xG�k��9|"<�YEZ}|��nZ*�n��(ٔM34x��3�z��R��M���dA�y��:��_r�d���}�~�Vg�t�W�V]�"���?tx�C�[J��[��LX8v}�1j?�hzbSԻ�	�}�����vb���״z�y�����E̼By�:3��7�\B���~���+n�N��B�}�gw���zeYCgɕ�[�_�p�]�ae�/���hIk�~&;�ǟO�<��1���he�0��r�X3�U�2P��,��n�d��`03��`�I������Au�4���L�'k�KL{|�>��a�$��6&٠�̄gP7t���{T8�ë=����=Q
�T��Ւ_�Z`pm���!�������v��/�
���?7��c��hh�1��^8=��?HƟ��ll�{��d��A+&	����؉��(,xx�	�R�ݾ{��r�MJ�cQ����_B�샶�ɷ�S,KgMۂ&@�ӏ/	8���&��/۟;"�r����E�E|1e����؆�bq����P�:�m���n?1��
�����3"�el����6I��5�a�M�C�pA��t9�%�7ߋX�&-j�K�����ðZe�9�mL*�뷖�z`P�xJXB�a����h�����r�;Jꂍ����n/�����gY|(�������O �jb�+}�8�݁��<D��.�@���`d����Fv����5 ��7���F��?\Z��"��W�
��>�o%� [��юN�Ӷ���@ȴ/׀��W2.�L���������6{w���^��{�B;I\>��C4>*>s�k��U���ꒋS�Ҟ@�iU��n�]�j3jq엂�95w�z����a�\ �P�۸<R�5ҾZ�~D����m�6u�E%F]�^yVŹ��s���	���2�I�j�[�z�p�i�U&Mb�O��;lCz��z�ޢ9���[ׯ5��߷�3K�8y�'	O�W�S	��^X甫}9N ,��ݺF�0�^�I� te��·÷��ø3�|���u-�MAGa�O@+���4�4�����:|`Ol�����w=�1�_��J�7�x[7��IK8VK�wH�:%�$�`�拹 ���5${���S�/)].F)���9xMX�hKY$v�� ��%�����`�~�����K8,�1�M,��[D�dW���e
/�-�1N��6�yL�9�Q��D�Y��B_	z�^6�I5lz�.��D�U�Zq���]K&+�����<�x�x\�P���+��l��a	���A:-e$[��|��8�<������IM��񫢇C&[��\���c�7ű�}M� J5�U�!2�Ym+2�X����[m��l["����� ��4��c���<ԥ����f��RP�i�x�"��u�'B����Q4?c��R�?%���bb�+��P&�2�QK<!�ך�ZX�����Q��K����q��!�f�ʑ�%֊!IQ�ճ���qd�C�u��ލ�C�47�I���eȩ�KwtW�T��i��x�w��}�7��3C��e�5b�Vsd𖃈���:^#Bw�ɿo$�hS���N�Q/�����%�S��R;۶�2b
U�`&.����n��c�}\:���$�Z�xL�3��ţc�L]���v6�o�v,�IC������3������Uu���<!�4��x���1�tv�[���t{�Z��Spڛ���S���#߁b�Q�3eaɎ��m���$j��=�K����Qg�Q�*���䈸�-H�Ӽ㚢�}x_�x^zC
���/��9��S��^rL��i���H���#�h�БX*����%�}��P�7Qw���&�a������A����\�fa��o_���Qc��D�A�{-�O���`Q�ܤ^<$w��|��'��z����/Ч�	Z.b��D�a����+<5��p(�gd?�T |����/C59謠����:1�/ �"`����s�tX��*dB�%���K�.1V���	��q�Y^���W�9�Ж
�/N�j��I�a/q�ؘc�d�u+����z��`��������&(�ꟑ����J(V^��V�<l%��@x���ў�	h8�N���E�4ܜԝ l�.�͡�(?�~��Ğ�6����ڍ�o�}J�S��J㲐ڸ/(���ﴼC�?��iF�y���:[�}�t|
�`.�S#�Z{�'�[L�����G��C�8Yy�n��}�F]��
|J�����,�-4�p��vM!H����=���Fb2��_��6�EšnwS�8}��d���Us^ Z��	{�5P)����m�S�=��}P�'�eY����㳴j@��������:QDF��8m&|�T��9R:�����l��^���E�Nz{���d������VxN������Ѭ�цkڞ @�9�B�we0��f�%��2��g@j�5��Q�Hߓ,".��VSF�8�ĺ��	0t�[<����B�)H1.�3�Q�	�U>)4��f�^B�m�<�~I�p����2��f#Ȇ�R���m�Xca�i��)u�O�@��)�,��KRF��K�/�� �D����r��Lo��՝�r�x��Y��Q���CUD[�8R\~ ��8nh+�T�/F�?��)�, >������ֆ�V���r�339�-�0Vŀ��q,�A��h�O;RT�v^u:Qt�!9��f{z������C�W���� �E��f�Ȁ���ox`���12�{-狿�6�G��R�5@�-��&]t��=�q�x�-e�Q}��n�Ѻ�9��X.,�QwY���ѻ�Ə���$��q0��������6��Y7p�
<�b	�~+F?���H�)���L�
owa��^:XYů��[����h����s��W�
IMJ��hMR�rc��ԁ������`N�����-Ƀ^U�]��y΂�oQ���f[�m�>0��e!?(0�<V��ܷ�Lta��{�#�W���4��)�I!}GT�jB��Z�4^�,��	
;r,�'�)R��?�5�����Vf�	 ���{���6�`Ī�`���睌&�K�hp��%K���D��y���$B��w� qN،�Og����uV���G�pGI�G�~G�PļT;-�V>�|;�eDJ���b Ōl?���=��uҫs���m�^�|�'i�j�+���f����3���17c�^�{�F����\pi r��	��s���1ܟ�_�{.�x��[����a)N�1�i����TĮ�CD���Y=�z#��/�z`o鹧��fG$3��y6�w���9~��\#1�)��;'�5�����	R[~5YH �Z�[ �{�@l{��}���G�FȖ��]��=�z1�qȬ��}��N���@��+�� �0�Ք����%�����i�E<ՔP�c����S� �!�X-Ra�:BVi!����J���n3��e0a���žb�b�N�4�a&G�"B� ����V��^2��}-kO��Kl�I��,o��#��k����V"'��Ud?{�P����>�&!.2��5�t4��o�t�܊�|�Z^i@���_̉�)��+͈9
�$���\�
Eey1�eʻFe$bW*��a�������O(R^�x����qX.���L�IaU}j�q�klM�6��&��
#P8}�~�W�5ĺ����(��t(�x��/г*Y��3h~m��Ɠ�X2������������wI1NS׿���Zb��%4߸�\V�y����V��r�Y�ZL��S�ᔴ��L)z.!��j���P�"�1)h���@�i���8�Z��3"U�:bG	����S$N�k�T2Go��.rP�3�`�e���bH�;	��z�Ԝ�FhHZ2���f����6�fq�C�DmFY��0���I�	�Ms��BtWvk*��q:�Z2'�ӐD_F/��"ѿ�lV���DqOԕ� g�R_��p�L��}&(�F���!���8�'��}�>�V<�M���V�꺇���P��)�o"1����}�s~���6�tZ�FY�:F��Q;
�@ȰK�.#a7�aC$��|�4��T/tb/0s3b�ZdP����W4�UCʒ�ηw^���{|�g��)��>�ʥ��exgK���v�;.�gy,n�䁪<!��
�-B��I�"-7���ی��B��:�*���[Ϳ�tT:(ôSu$w,+NT��|�;�r�S���`��D�oH$W��+�7gұȯ���Vq�N��<D]A)�l5�8p��e�9=i_?r������;���Yo�)��	�f��~��jT�ܟ�Q�O�s�󾄀	����������~��x����П�����{��F��H�����)B�w�6g�(RmߖFg[J�ָ͞ݹ/���Z� �.�������lK�}������5;�'�kd��3���A��.?:����	�$���*|��F�lXv�.{xB��!�>'�$d�b;o໕>��a�7��>�M��&�/h�����q@wr����q�țO�4yg0 ��2΅P�f�Q�ټc�/yr��Ѷ8�H݂u��|�P���	Z�ѷw�Q�Q
i�b�DJ�B�g��)FB���SXh��l��o��K�'��]t��=���xLx9��'/ME\ �'�atx���Y��-:1DUD<7p��3�c//�VĒmz$��5�xn;P0��l�DtR8A8�ۦEܙr��Û����)��x� �zy�>h(�e�W(F��zy6`&^�C�iYu,�pP��*�H��U��?Y�$�g�\�/#<\��V�q�@}�z�{�s7����A\p�		h�1'�24ϖ��߽;;d|V���}�J>�T��'J aQ���-�,�N��'e��kc{���Q�;�U�=��PN ro�<6�*y�@����J��Z N<���T$�J;�;E"J��)� d��4=}*���,|��H^�"�k�o_A��cR��=�����ebs}/^�z�ŏ����2
	�.��}Ȍ�@�J� ��	��玖���=��d}K%$���Et�&3Gu7r�=g�>$�)Ӊ�l� r�TvM���6�K�[Ԡq�c��bK�u� }1����2ա$wa�����⣭Q��l����S��SD�=g5�	�)���䔵LmԀ�/���ZV��ݭ;�ta?�]�2w�0�
����ة��	~�;5�N� 7k�8��/�e�o�q�	��.4����q�`x����������w!q�j�{8<����.�/�U�q�Z���,i���Y{�z>P�E�Ho�6��W�r)���I,�L#t�j��A�Կ$�kz���fX Ī��5�[�Oy!.GN��N_I;�X��x񪗶̞�n�^�|��\��m�GS ��x���2n���pÙΠΘ��}�4.RTM��O�%��R<ec,Dt~ې�j��gi��^���B���y�v\��d)�q�9�Q�>�𜏙�ֿ�ߜ���h�O�g�g�/3I��Z{dI��3�@�=�9��u���'Kh�<�ب��s���VX���Hh�5����Ql���b��0���)7O`؄�%�t%��p�QH{���7I�a��%�@���i��PZR����Vռ�&�����bC�*̘Ԛ�e����F{��L�b�W�^jV3�W"����PE�>���`� ���O�c\��V��˟w���usl�r/�#�Q�۬���u����Z��BN�.�r�6'Q!���3��i��%���Zy{5���u3R8��5	���0��hԆUƋ�Lw�Rg�R�)�;�W`;�G ��@�7*�bh!�����"�}'ϯ* ��^>% )w,�C�~�?6�v��ԥ�n`b��F�]��8�����tt��]�Io��cR����L���[-`G7��)��N��!D��0U[��f/8��k)h���T�R_Z���8V��ف\��ܔ#�(sӂ#���w�N�ld
?�~�G8A�mr��w���$��'��N�;��G��F��~�Ñy��ٗ6J_m��]&��������k��Т=��W��G�˼Sqo4^}��x�����*�j_�3o��|X�a/E��]>m�?k3��LH�`��\׀�\��ճ݇�Z�".�9<u0�Ճ�Q�P���j_ ��I��s�����E'ᵌ~���F��f�;���0ӱ�~P1v�ߍ��J־ 6X�M��Uaԅ��(=��N���ZV�<��s��6����	�{�9&����LG�&��# ^�x�Υ����ü�8�x� �=�e��w	�SZ	�3\V�LN}E�A����e�.�k���S<s�;:�c縬nz+vX,#�%O�@$}dQHL�E�@	�K7��y�Y�M�!R����4>������'�j�*��^�MiVb��t��=��U�H��;�y���
��("م+�϶��K��Y���	9 ��/�n^Ek��������u�13(���|�KY���~Y"��<�c5a*5j���"�(`n�H����r���iT[9|f�d<�}8��Pwsm��}`^���|�D���y/D#�ߪ�3K/�-l,!��S���r6�?�O_Z���@|����`�K���a`&q��mH��'�8����l�VdoD� ��kS�����*���c��;��8����dE��:ۮ�	M��]�~*.��b'4��A�(y��|�z�B�1��9QO4�����,8{G!�͞�o��Z<!�aK ���H�2�/
b�Y���pKG����*�/�1!���UB��@ ��L�|��N%,6).A��MG�*6���Hɱ>�bTBm2#%�˲��w��&eɺk>ͪ:���nd�ITҵ����O�vy���^�0�*��$��.!�9�m,]	�9 ���BsXu�f�L���<Mm�2�!	N{C�x=�K&+�B�&�%*��'���pe`�}������?��U�M��w��5���h�대��R���P��%vX���]��$'�-��Y�7��➽�	�����Z���5�a�@
�Őd ���t����h��No����6V�o �=I�����E{�-���-d��,� M���(�o��Z��4��[&�������0%L�g2��?hg��{���/�[E�ԲY'��"�l)�rW��FI�<�����&A����P��Q��.�bԯ��	��p�٨+��-�ӊ���S�ϊ��ϕth�C�4���Ze�ևl�hC��qvm*T4<=���H�'7'ӣ��$�~������coj�ˏ[�ΗMMJA�u�S ��Y�KC���E���q�iaOy[�ZM�Y�VP�d��ѵHnI�`���q������$*}�]��IZ�`Z����a�I慗w��gW��& ���nS��6��|ۥ�<���X>�Q�*p D�}�沭kx�\��F-���k-
���e���4���|����-���^U��:�N�ڝ���I��`�"sᰳ���?�F��a���T�3.LIW�`_L~�q]�Oo�.n�2Kyb���rB�#B.5H$�霒�ؕ���m$�Չ�w��U)��vbw���}!�X���Z�S|"�~�ͧ�@��/}'$�ga������;I�A����u���/�tE���ӺA��w��pS<�������mJ��2�����W�;'�H�U�-��O6b~���Y��q�ۜ��A����g�J9{�n�B�J�KrZ�I֮�8,��%<@����������￐$ɣ��5�SC�1_ue�"3P�N��`�g^��H�<*�� T��E���P+�xl�X>Yȱ��g��T&n=�Q�����H�Dѳ85FuV9��~�[q+/�F�����$���.ʥ�i8v�I����j�ǫz����'�="JpU�w�1=��TlV�s}�K���2�����L�<D}p��]��8I�V�N��t�6�'5ɜ�4w��X��+S��|��36r�����WKg����x����Xj�� ��w ԥ&�工k�vOn��J�|*��v��b��)��~Wi�W�ՙ�+EVQD��6��V�F�Π��587�n��c�]��k�z��1E$�A)H�-�O� E)�C���7��w^�^��^��~����sv�Q�kh��ج@v�W�Ix�H}E�,Xͽ�_h�V��XYP`��8.|��CVjkO�q��C��+ڍ�oJ*^OH�I��`���VF^F���ao?���*WodL� Lzf^���V�n�^�$6G���wyߖ��l׭�)�������l�����o@q�e^OEh!����[��&������QQƪ��$9㡘-:�X�%Nr ��
+���B���K l V�B�E��XO.RM�_B�d�p1�e����h�Z�y�S#�@�u�Yg�?�� Ca�h�L2���f�r�:�Bn���PCx��ͥP7J��}�B"��Q��0���V��ծ�q3 ��ZWʈ�����x��3c9~�A ��祲3�)a?����U�G�s˫��C�BTe��I��m��ʕMd�|/7�W�2��[i�<���Ɂ2έy
�P�)A5��x�Z�5�J�������SbT�W��HL����߭V}��S��ʷ%�8Z��6�;���U�/�6鐒_j�/ף����tl�j��\�S���$-0I@0��tw��m`p&n����&V4wkWsæ!������_�����e۫Jy=n�g�&*{��B��hWW�3eYʸ.g~��0	~ț%I�5��N���@;��n`>0�3�i��}Mb�	�f�x�]�O���T���ɜ>	!f��wj�vH�簚OR�IWw	��J��g�-Dx qs�|!�Lx$\�}�C-b!Q�n��%�Yr���(\t�y~4�$�`왖8o�4moJ���l��&��	X����i�����"��yH��x�R��Gi�Ws�5�e�;�s��P�R|�^xt�O��G9�(�������ٕ���X���';2ۈ�?�ڪA
�1�>?�a>�,��z�����2"n{��(�'R�"���KtcJիr��c|����z$��O������V�s�*ZYl�����2�XQڗH��D�*ax��LCO�!��~���ۇ�&��� _>d!s���k{j5�ą��u��f�/!�/�����0z<_�R"ߌG%�a6�ȶ�Z��!�tG�a�ԫ+}Nt�4x"�arq�5��'y��=�R^Ѱ!���p�bX�#X�T��c�G�T
���l�U2���r��M!�7����ܜ�V���,�6��8�Ʈ} M )�v�k�3Y!V�Ľ�<��� M7M�I�TLovIP��;>�s��Kalƿ��<��K3������AbU�^��[(k���MՀ黮�ls8���_[c���5�C�#B�8��������``Q�m��>>%yf�X�D V~��X'V┋u}TX7(���}�#&���rϾrjryLL�Xy��a~�M�4r��2��� �M��V>lt�����z�Ew#� D+?��9K�n�ɽ<�k�p����ѵ��ٟ#@xv�F��vf�xk�����Î#s47jaۓ[�פq�Q����[�$1~�.FΓ��-b���Ap�������g����'��f�z4>��N�{n_���k�&��tF&s_���'ɒ��zE�5���k������7��5V�&�B��^�0�\��QҰ�/G����o�k)��4mEѲ]?U�Z	ԘW(�}�'���R�;���ǌ@K��Ϳ�)�/��	���i�S��B���4��X�9�]@��YNA$�k�7�ۄ_�*�8^x��7��}0���2G0�`�}��8�У8��hE�9��;HT
���V�t�cV%�;1�{ձ��?@�&�V����(���>2��MZu��g'm�U�P�(�=���0�y˷�k_J���*@�{��ٚ��;�j��q�D�W߭���#8p�V2;�̽����,��7f��d�Q�]������ZA{-m���:�dM�x^nU��H� �G����:�ǹ\��Lz����Ò��bu3&��J翕�Y��٘s�S����#��Y�w�5��n�X���?YB:
�����׿"˥Z����֗q&I�/��R\�`9]��˩e\��ˡ��ׯD!P����z#A{QYsK.J��E�MΘ��+�!�0lV�@}vǶġ�I�s���Nn^k�7�1X�Q��f���L;w2�`qiLw���f�`ϚY�н8�9�C��WΝ�(p����?b2�������q�K8�:a��Y�-��\Pˍ�-m��H�z��s3���%k��|���N���/�%���# ���]�����4� kޥU:H|�,�HN�"�2��.7H�y��%N� W���D��lR>=-d-A�E���`�^ ��d��C(:�k�l�8�e$h�w�~��"ٔ$��/o�Mo'S����e��e_6����GKҶ�d�ge�y��D�Pջ�O5`���فy"'�'�����{?U���jw�" !H���A�;���Q��feajZ�z޲5�EBG�¶t4&"���������V[Cz|9���d ,P�D��4��?aCѾ�E�R@�`�V�y�K������Z���J�9��x��V\í�LW���2��'�k®�\Tz��>8�jN!��7�����!�A��+��5
ŝ�a
��p7d���Wd�T�oN�Vw�ֶW��7�4\k�y[�1w�#�N���D���^B����h�yR����ǜ8,�
\�^ +yK~қ@� uV�~�����vZ�,~T����J�<�KL��XFR\0�B���f��`�K�v�袁b�ܔ5�bŽb���L�2�.����Z)W�'n��H�[�Bm�����]v[�.W�$)��[=Ԍ0O�AG�k���Ð3!U={n߅���?T�@;ϠV�@���e�����j��J�?B�{�<޼^^����f��׷���O�t�O)5��怌�\;���C�hЮU����>�(��ǎ�?pHd�nBt�!�D|
���d�H� N�-��k�=�$Zur�!/���!�,/�q�e�����Y0��A}��2�ۼ�0���6��}1ܧV�����-R�g䘍K"��R�X�|�W��|�{��M�R�X'&�%���yX-���%��Y�}l3�$��h>�h�%_�P�3�?}�3�5���,�� �R^�����/��F/���C�$<��A�bs�`lH�N�I����yT���qdZ��q7�L�"y���"7��$���_��p�䈩[��#�Ǐ�V�C��}"�G̓c]FeW#�*�%W&����M�(n`b�Vҕ�f|�����H~����թ>o)�iL���%Lߞ�	�~���?y�W�é��k�Dr�E��I��
f��e���u�q�H�-��
��~�gJE 3�Z\��n-�i�oŧ�d������aS���L�&���U���5P�;t�t�[������]���T�x6��+��5ݘ�C��w~$�$�!���bv׶Ƞ��x:����;z�Z�D/N��"C,�ܿؼ���g`$�e�S˥�`���"n�S�Ub����%���u!,�3d��0��R��3�=�^Lۍ$��nl'�d�C�
5|��p�z^������t
�|bmU������<�e�m�~!m��YO���ry���׍4��cc-��P�.'E0�t e��-�T�'����w���oZ>��d����d�r�x��a��Q�^��K.<F�6P��7���kJC�o�&�X
u�}TO-��SyN���#1F�f�"E����Z|4�Cɢ�kX?1Eҡ;J����ui�Ȍ�,��5���,�G�W��Vʱr� �x�oP��'3����2i�[L'��,�����
�5V���|S,|_0[�ttm�wk�v��gG�a>�x��TP��L���GlDȒ�^���}���ӈ�� m�T���g.qJsy��X|p�'pM�n���x�RO�G`e�4Yv��e@C��gWz��t��!y�>/P���4 ���Ȏ+��,:�<�D i�=����z���o�?^�`����Id�8¼3
���[�4�b]�ш7x(�ܦ��5�x`&�@��>͞�gMMM�-j�YAͿ:[FV�|��	��5�v+���Ê�`'�5wa2��F�Y��N�@�t̬d}c��i�Fp��)���'��XQ�6M��~�5��"�i�7���ͬ^Awy:�B�ϖx��Teb�:����dJ�>������s���/�߱;o#��u�t���WD[-!��67#`G8� ���X|�b��լ�)�l�`�\����A=0bOI$��[���5���.��ն���
�:����?h:��0,�i�����l��d����x�J�̀�2'����H{;"�c��]�٪;�꬐�����o\���}͕��wX)^�m�ljD���B=>��gu<*���e0ԝ-�n���s�oo��6J�;M�,(t��F�T�����'#&�ums.�LO�%R?�Y���(_ ��5ai�4N#��2��:�"��w��q2���-76w��;�~[�_�	JZ�7��l�]m��b����D��� U/������\Ƙ˨�j0�g����sb^����ʲ0uC ��	�d	�����x� ��+[4�׎����:9%��$#�X	��}R�ݺ�p�~]����pr�ʙ.����@^
�uYZ꧖�L�����q�����l�V,�Fg�����ef�8�Ej�>A�,�>UI,�.��-K� *��y��a.}����Z�3�������w�>���s}�4n�l3�@�#�y^vX���Q��>��	y5Ly4oDʷ��6j8�q#L�6?�W��(�ec��k�G��[L� �ٝ���ߝ�-?$��آF�IJR�x�6E�chr������$�>�3����)IQ��+J����&��q�!<lw�1:XVxC����u�]�;�/�4<|��%Lݦt�g�t�Eb��P������Ls�1ڻ��ݭ�5���9�~��E��?D'k/9�ѩ]ek�&a�X�����b�Ҏ�����e�p�-'Ie=y�m��u,u������/P�݈��b�v?�jø��T����øz+�_��D2x�i-�V��ӂ=�	Y&сnK$X�o�L�I0r6m��P�qoHy�l�әÄ�+�l����X1�Ӣ�;0{^����"u�<� �HW�(Yz㋅�s�?$'�^�A�u���f�bj���%o��8�Ũ��l��%��AI/��H�h^�H��{��w�. �R��Ю�Oh
n�/���
�%�r�;�.��x��f��,4DU4��cʬ?�� �M�ؘ��i|gr�
�o��G��'Vь�\��1]Biʰ(��~^6����8 ��>��~����?,�ݽ A����kz�&t����/&!��E5�^I�XA��R��r�}���%�u�v�-��E4BT�b�\����A�
*3��^�T��gC�JA~���]S��t�9,%��uI�;ҳ ��X�܊A�D�E�L ���h���h�R���`��Ճ��%�Mga ��QXU�|�qd�!�E/%��i�zcl����>�%�����X\��-Ȯ:*V���Y}B.X���M�����������8:�m���KP�2�m�C���Q�j��\�
T]�w������L��I�+H��7I����s��3I\f��P.⋃���,���\Z���JO��>6��YX/�̐L�n�@.q�4;4����v���E�O
�db״u�H�{7�.%�gݠي���X�S��B��Zc�ճO���z�2�2'���H�0U4��
�a�P�	��,���O^),��,����)�,���%f~
�q��N��A��`C��+5��I:i�A&��i���bUk�4D��4p�������ᑒ��i}H�(��O�J�s*���|~�+ć�C�*�stI�_?�c�q�����6בX��c�����c 	�Y���Cב�(9R�w��r��"¦��qU֋��xL�=wȫ3�:mL�U�������Eʡ��V��P��4��sO�,9,R*�>�i�W��MGz-�{�N������nzG�z�9�^O*���O��dg�7��s3����q-�-O�s��;�L�7�=c�e'��GR��'�|A*��ֺ��{L�)"U�Jo=O����~l�V�R�]VO�C�E���yP�}�޷��W�$����=wa e-㘐�������g,"@㺋/��s�(�E7�>c�\Q�e��2h3�z�x{�1}�;SR��J�bCTBd�q.s��#Q�ְ]K���\���z}��x�Mc��҉�K;fr��}>�6\w�B?�&?P�>�D���g��su|��ć�z�/������޳��.�SkC�)\��ltƕ�/sX��(�IY+/�m�XXޒ$�<C�	��@����U��GKJ�T����P޳^��;z�����5��"rϔ0xGۻ'��\L�f7������k����@���<��Ͱ�g@C�nA_�O�� �MI,�be�g ��*�~w)`���=$�%񕐴�ܷ,��0��eW��̤C�rD��=��b�_��̈́z-�'%�D��t�!��#���t��l0�M�`�΁7 E9��c����xkVߎ��F%o/��H��O)��վg��5w��ή%��+hh�����#'Z�1�P�U���!1��<ט�<|x^��&���Z�>6�̩�������3=���ҫ�4{�rz�e��T���M?��v��D�d�5�od�=-bh�_7,�\7����dun��x��ے_1�k!�^`�BD>�%zCL��W��H>KR��U��T��e����"����m?�ϡ/_zV-�e�6��>N�DCj�� �)L�k&�뢙�A��_ON��7�21`�f�Wќ�O<G�����t+���:�3�H>	��};0���@�[2p���F^��»��@#��٥��`�>L;����?��8��fk 4�$pך���a�ʵLm������@�n� �C:�D�mr���ɜ̡��LZ�ۍ�$O�[ܹ ���/��мYh1���6��Hf��^��B:�f-ҙX���B�x�wx�;��#��g�ؒ<�U&A������M%�nԠ�:3��Ӻ�2o[7P���эh8����r��V�d4Ѓۯ�Ԝ{\��u<�ao72l�5�6_�ϪD%����M�}#��`�%�L�s~4�5��A`B#X������?+��0@���=$�,���N�$�H���eY�j����?�W9}�J7���K?�ܼ�	s\����@�:��,���\�f�	�C�Y�	�}��=�b�	���\�7~|�1��F�6B�F�f�[���qOЬ@��(k>��
�ݖD]��.�p�'�j�9]��5XG��ai��F��R�;�U�Q�oy_���*��4�]6�oCQJ�~JCt5=�tP5����Z�T���A���'�P�v0�Gjv[U�������7�)������f;G�m!ɦY�:_�����_�k����N�X����1�FU_�/3C�GL��)'�����)a>�'vC�3;�hN����7H�P��J���,
v,r�p�`E;�l����ԇNZ#����Tqa�����II��J�p����t
���H��^W��cyAt ��������(���������D�e�CV��E��Y��/�to�q��qS^j��	�+R�f�`�ܻ8@r<qg�L�=t��<���_�t�F?J���
`>���d$մ��O�ğڣ�~�14�~u�2c� ���u��6,���
~wʏ�:��x�� wd?�%�|1]ļ��ܶF��)�Vf��J����a2ԠTe�W �]2W:Hi�Q��,\��X�j��w�R�B�/�u�H�Ҥ�u\�[C�B��_��d�G&{}�ƊHZ ��L�PIU�^�8����������d��#�F��el��"����e,z�w��^�/86 ��ʃ���9��yJo���~��#2gth(�gM���3��K7��T��L�d��!4�b	z'�"���hL�y�?w�,����SL��|?6�%��:���齨 �3�\���	1c�h��"
�t�1^[��ZQR���Mv�֭��#�tE��� ?���=��\d#d����gV�%��H�`�����g،�(_�Ȥ���m��f�P����59E�4n���=�<|��]��|I��Ibx�{f�*Ҫ��v��yS�I>/��JiE�B��x���X�0׹��'QT�R��I����y�����9u,�W'�|p|'#�{H�;n�R����$��|Hd	K��gC�I�J���'�T�N��瓒�\��I�1Z.�MT��=���k�nZ�C46ї�x� &R��F�������.�1
-�sW1-�z�E�w���ӟ���m�J�Z'��y1U21=c�.oI�g��%��sL���ul��*�py��=�c)��Ǿ�w�f���t�����t��6��	%]1K�߲��&�s��}�A�O=61�>�SD�c
������$l�q^�ѽC���~/?x:��>���j����qwj� *�\�xm�+��]�}�Y�N4JH�|Vps-8%3\-��?��}W���Zb��؏�2?�_-�0L�K>�	_���l ����&8\�j����o�b����Ni{��	��[x�b�C�-Ӌ]N��f�����0���%�0o��=(6F�$�>YQ��y�Ui��l	��QD�Z:�JƗ���(���L$cG�`����(�(�Wu+5�+��sg����qtG��!�����S�(�Dh��E��/X��I��
�PȰ�'�.I��P�h����/�h�{��y��HS(j:���`��^s7�������F�݃�$�""��39ɡ�Ig"���V�&���M"S@������<T�E���6��<}�fJ�O�1-�wI�J&@}L�WU���<f�ַ,lgdbLH�'0��Ac�4a������5%�Fl��ە��yi�l���0���z�Z�c�&��M ey�{*@w�@���	r Lz3��X�$p�=�1�� ��QyG�)Cʾ�jP��YMG͸<�����Bs�D!D�� h��X:��go�X�����kbL0�Q`�q��>�ty����"���5�R�Am�M�sX�
���&���^�j.�e[G��^�O�n��%�Ar�^א����y�o��J�ZT��Z���O�*b|�*un���,����r5�����a���2#�S���Nr�+�̸=.�hSd3���f�|���r�G���䄲�e����!��V����r���@'I�y�=0�۰8œ��3w�T�`��"L�8�B��`�\S-�[!g���*<D����W�U	�گ��Vŉk3b��(���`�}Or�'�ֲg�D���Y3���^�\N
%i���D��&�fKS��w�0Փ��.�~K<�q,|r��M����,���kռi5&p`}�_.���t9~p�s�_����ϊ����5��A��o�=�1��>�*���k��R ���<t�y�7N�ÿU4�I9 >�U%�Ie�%ޑy,�מ|�C��ċ�����K���XUs$���4���_40��W2�Dd���L���9FN#�����e��k���L]�궄�9yL.pGe�(��np'��_��n��킓A�F�����ɗ��p� J��Y-���Ƅ�t�TX�HQ"O��,�t�:ٛx�сn�����Bc�҈F�:���8����y�_��CZk��T����I/(���Q%Q��=:�B��	r��I0�4�I�irXt�r�W�H�r�	���{Wrȧ�4���ta��W~��RQ,bIHJ#�i؁�`��D�ͱ�K�2#��4����9��K�̥�#J�%������"��b#ϳ���yh��)�%�p�,rfCf'�q�Q�pM���,l�+#r��h�CԧG�)��+����1H����<��q�,�|�f�Y�C{��� �����D����}X)�ʁa֜{�����ԉ���.��Z3���q:Б�)Ǣa�|խ�5�{~"o�Hr��Qu�y��/}����<q���ՃrϦV�uQ��v�N�!��xt`ڮ��!����wV���8�2"�B�4�����"�r~c��R0�cr���!?R�\afl�?ب�"�̕���F�oi_���2��x�R�6*��(���%�����*���}+�[���K�`x�������%�f%��1W��f�Ǭa�2�l�gyZP�����!T�� �e��1>�>�K���U�1�ݳ�*_�5�C�z�:���m�� ��?9��6F;IfY�̉�Z������0��K�S����&Q,�@��UqѝJ#��9?X�ۏW|0P����~T Q�\�_'TGJ�e����Q�5�����&$:�C��ò�_7.ZWrcVN���r4�,P����fԛa|Ț��[�:�caAjz�%g����:F��������m.r�T@i?��~��8�M'����3%$�#R]]D]a�ƅ§�+-jA�*Q�o|���Nq�A#벧/ݏ�T�	}�T(]�wr��w��W�؏��zP�>�m��ܾ9*���R;u.~8_�m*K��>�����-�ﺘ*J�BW�N�i`^f8~mw>���>=i�6�,g ��\lT��R�V�����[m>(�*�j�"7Oz/�"���K�ehа���!w�t����iw��D :r��GK8-����P��h�����(tS_�j��O���qh�+)xf�흊�w�L�b
�_��s��k��+B�����&��;�5�C[��D�=5$�ǛxHI@��f�#����oJ
�G�q���Nh���'G+B5��^���TF�dN'�����Ӄ���.˜9�%N�/	-|ڭ�r>G��'�D���ji�}Q
�`Լ��vm����t���`}Q�s��/c^G��jm�X����@`.�z��H�!� D�x#I*� q�aފ$_˨�����b�A��%��;݁ӴЛ����½fJ������̧�
/�({S8��;B��DXekg]�N`�*�W�U�D��g���S0Qy�y'ۻ���2��7�p�)�#M]�`�{Ư���D����KD��>[>�"�2�C����Ul�K�pR��#����J�}�Ҁ>�Z���!��{A�|X���sm�f)ƒ�|j�!��S���I��\�����B�N��f*hn��Ev'�|��"��%E�Rq ���$1���6����QZ�Di	��y��p�z���E�����[H8 �:vLw�]�V�	�P��1���=	�Җ���F�G�]�#�(�?-~Ϝf�b������A���+j�9J��Atr�[p�B��{�Sޭz�~�˞��?`}׺������E�v2���l~�V��M�	 �lN��d�� b�s�%H�=�� ��-X�ΜHa@���섨���_M���[5�!�>���aT���-	=�w�vӽ��C��?L��%A���e)C�-N��pv���+Ί���3"���ب.9�ZlS�Nㆢ����ڌt�t �Ϲy>!f��{�U"> /w�����i����"P�C ��W��`���H�Y��N�8��a[M��7�M���Dͫ���4#�		�1�#�Zu�XL{��Y�Q�?�QvFS7OeZa0�	�ޘ����px�(�����B��5��`󰄒1�{�V#9A4|C���g�����[t~N\� j��Kl3�E�q�{�Vu��I΃I��HY��]���^S�M�e� ������*�V>Y��r�S���߳k�H^,^�n�?8�T:�p�����h0xƗ���M�A�?g?�,���'L0;/?��=	�>�{��.���W&D)L��.:դn��u9�|�خv�Tx�S�{�������Ƴ�R#�yB�pq@Ʒ]f���Cu�:�	a5Z�����A�f!����P��M�)�;!P��&?��S/�:�}D�)/:�s��AP���(�B����	#:v�1Z��]�kX�¢=�nLb��K�[tk���i�E:�������5�.����p�W[@�x�����ݿ�;�qd5%배[���4$����'��L�Ӵ���N��V6��'��IyYG�bj��~&Sv܇�LN���pK.�Vw�X4-�4�*����kT���uUf��zl���F0��7��R\����c~@��T�s���2�ۙ=ctG�G
G&���Їw3ႉp*�v� �1��k-�x�����PM��?��iT�̵s��z�ʥ�DhD��1��qR��U���� ���)\�����p��H���'f��M�+}�(���J��]�-��a���59 ͜����!�%&�|eš.�W�[�aְk�u�%�T�d�*��t�bt�V��o���g�!%�K��;�p1
��-S
�.b����C]N�J�eۑ��d��f :�:�M���W;�f$E׍v�ʫY���YνY�y�/9���2�_����v�>m��������q�_�>Ś�V�Ӯ�Ǽ׉����gǤl7T�T�۷R����τ�9Ґn)緄��ԉ��Q�f�ۡ�{��߼5�P#�9
Z(wX���_L�"T���J��[@4�,�}p��*��e�wT|�Ŝ���X�V`����K�z���=K���K�6�yJ�g���1�����\��J_���#)� F�D��
�l(P����g/����;�2�Qg~{���ym�p3��v��5NOD�")щR�S/���}��ǐV/f�|�k��C#�3�������z���1^w��u����9��yEe�k(���qK�iWw�>: I�1�FVs�\o%^(\O�f��/,h�z0�;�R��?�`�J�;��1(��-k�;�����3�d:&-��u}��|@rQ��t�P^�$�I�]�B�Il�C�-o.#jz�F��x���#A��`CY�,I�쫮��r��q����H^���דp����wL�� �+ (���g��5+��p�?���Py4XǴ�p��`�{��I" ��na@���,���Y�V�JV����=������$j����`�p,�)3�6�޲٦J\?�*�\���M���BO�:���:zgY��O�ǘW�ju�Vk/���]�Bi�֥k�+ij$˻� ��#��G[�߇�/��h��΄y֎/�5�ꄉ��>.a�6q<tBVK���NS��>r�Ϥ\����wl�j��)̂��4������Q���%�_ļIe�j=ϩ?8`{�
�k�Sڒ��D�>X�˻��8IVw`�L#����x�`Js��b�ʗ��R�Y�M�+5�sש̀#����S��]c�0��D6� ���+�	k̞��o���z���j&��Z���
��۽�w�����-MG�]B۪��(���m
&��7ѥ(0I����rR��dAp�l��@va�toB'�^U }�t��ϛl Wb�h�_�o�0� %����(oN���1��-��*�%9M�(
��8�ӱVz���G~&��u�,���B��$]RÕ'o�O�	{�����|%�%�������G��R�����'�ZP�A-�e�<6��,R��3����{XD$�6�Ӻ�r�)^������;u�߳����a�;�#y���C�q������/�J��~�Ɋ[I, �y�t'T�hc���NH\u({#+xb!b�]I��BIXy�|6�E��81�:�B6��u�� R�c|�5@!�j��XI�J����#��Y��9[%�ޯ�����	\����G|?����!��[�L�+;�� �cG#��'�{�^`����炯vM94lbH���>Ƈ����:�`|5%�1���">�ο!���<�F�|��C���D�p�/)+_-��v���r���4��x�l�}WϹs�������	P��0'�X�A|��7�.�L$+�|�U;�'��\u�����:��u��bB�9�D H�u�0�:��'D���"uj�KwZ��u<dr�&J����t��\��Mê�C�@����	��6�PD7h�t��
l�5���i1�נNu�g�^i��]�bQ(��cIHt����6b��h��=)-~Ě�<�}-�z��L3�6����f^���}4��ҽ�+�q�8+�c��˥��Xt��nx��+�,X���"b`������H�>|H�I��ʀ��k���L���v[�h�ax�$�{� r_�;ഢ9���lc�G��[��W%���2����xg���1I|�A�qPp�o�|.	-��,&`��C��p"_�ީ�C�oin�����^��O�G9BUV�Z�3��r�o�-t��j�s�H�K������
<őv���P��pzǘ���"����#Q.�˯��U�S(h�?A㩙��T��K�R|`�|����w��?�Ż١�x��k�o�W�~�K2e����*� nQ�OGm������첰C
'r�}^�cb�xj)X׷�Z=�D\�U�9��/>���#�K��}�`,�?����t2�W�󱀯��=�����$��.�\�! �h-��qT�Vs�7v��?�.?�Bd�����3ns���>��|'g}�N���E�;�:`���@5 �Ǣ���zii�|�n���b484���3!A�bQױ�IX�ղ�]#�t&���rA��G��*��D9��f�Z��Ӆ��Hl˄)Yl�G�}� ]��F�v��á\u~@O'"�j�xh����T��U���n��[��*+55����?>�!��$'�#���h{eWѧ�Z3O����f�0j>N��"���1���vt�{q:��.X��W���o�
��s�F1
}k^ ��v�z�}[�O��ͤ��`�'[�Y�,�{pЦ�I��7���[�j�|5�h��>�-�9'
-;[�M�jg*�2�`�1�n=�ᩩ�U4J���ۿw����JcT2���kQu�ԛ���!�HN��g��-� ekkb�"���� 
�Ϛ�\��]4���N!b����+�A>_�4�*��=��?M�����D����L���yP��鈤�(�aV��nV>Ѵ>�s|0/Z���3{�S���`2�R`[q�7Z�'ݦ�wk(��k{*�t�|P�>��55���/��~�4br�u�*�`"�ق IJ���#��.}��^i����*�!���1�]j�	�Nh��G�M\�]�ڬ���̓��b|��(�t�=m�%��GseX�)�b^Ni<���{U��ڡ!�N}?��yE 5ȣ���[�GF�|w4��˿�I�����eG����>�>|��=�%=�1v6�;�3.r攤�*X,�Z��=9M`㡻��y�j���0��sɃx|P� 12y��A��_���vZV�jIȀ�ly�u����S� �WȰ���#esSa��%��'mT���b7%���M�gM�<г�w�uN[:؂�)F:*8~I����c�<I��u3ɵ�M�	����f����G�ڜ4d�v��\�n���5"�d;"�G��Tb)h��������n�W	�-��B o�k^nxA��Eu�Bw"�2G�W���/2c�ώ �F��\�5Y�QdK��nN�}$��{�wS�Vm�gB�}MXR} ���>�*�ջ�����pKD��&�x:[�8���sd-_��p�c��1�\V8R�}:������	2h�@��zu����9�.�]@5�`�m����T����/�j�|�K�uU
������=%����4J݉du���?:�h;��8�^���@�7��`%U�o"�pb����'��o�T���
�;��U(�'ݟ4e�����eBV.$��O��S����zD]w5�[T��n��^������t�>H�xd~w�
�A�{s7f+�4(�����M��1��VҬ�^��2���\U��]wG��.$�Ǡ�1M��I@�NK�����-i���Uh��-�S"�Х֝��(L�Dv���X�%Q���-߰>��M��^Nw�k�]������y\�k��[�5Rh���X*�)/����A=
�CГ
r�C|�K+0��0�_�4+-{�XR��F���/*Q�#�-$�/��e�*mM�-SɜMXī�h�4��&�F�Ṃx� ~���R��U�C�v���H��1�w�����:_����b���Z�{�2��w�F	${d��<���o����Va�@"w�H��_�
���(o������Ј+��_31�=뵌�6ۮ�m���T�/+����F��RX�#����F�\����l�S2u#��9L'�g�1 T�/g����Z�àQK~�Vc�e�[8����؄
�3���]]�sG��'%������o
�ź㠎`��X�F�-� ��¦u�h�V{&J9�4=�z~�XF��tC��]�[�d�ec��kt҉�8���A�\�K�v�/�`�eC��p3��rC�P'�)IS��s��1����:C�_<G�t�g���9����&�kf�9�`c�R�X�3��I��HO���YT���~��������b`��t��xٱ�x��0�b�v�����'����Hh�ɻ�풊k�|�B"��u�����|�"�|�k	�a^�L\$J��%�5�;0qV�M�!t�@�KSf_�^�n@un��CV��,�'�]��ّ�N��{�*bX=��{P8_K~SzhJ(>�q=�૎�6s/u�;���Qc׌��x����p}�f(R��}�u|����I�������c}�˯٩��D %F��7-�rާ�L<Jz�5,I��G��%b��v�p�a�R��wP�5��������V�
L���}Q��A��s�]
��5�}�ٹ�]�_���
i*�f"�l�^-�������\����r8����Y!O;�[y���pljZ�X�h����/�����{!�,/+���z,�n����=���{r:��԰��\L�YK�~3�|&U����L�2jZh�߼UBc]�ۖTfݒ0.F���	�-�Z_w�A��ԉ�ߥ���2�g����I�%q�����~!?m��.8�a�2*�'�8d�Z)��x��ϊ��t?�{뎨�ƌLDl��8#�:ǒ�N.���|G���Y��oP�=�8;��(ҨT�И#���,;xŉ`�^�m�^��u��C73P*0�����jT�WM'^�qQ�^�_8οI��zД=4&��#��9�,n�}j�X�	�ߚ3V��� nG��D)�R51
2�s ��pS=K5x�CQ;+?�}>۝DkϿ�w,�,g���T`7e�0�F��8�]I(�t0k�r�/	��K��
8"�aE��=ԙ]�l��4q�g��έ���ڼ����jsnH��s3a�g-Cg����j}.;'�c�z�����#�����#jxz���-;�v�6xU��Ph��C��+�]c[7v�������m\�dR;p�%r�k��M6j)
D]�4��p�X�7UHWx�#Yf����O�?ǆ����Q���g齇�����\���,�1���
>A�SD�㭛�#��P����JHh����������␜�"ۦ�+-��l"g����׺��vU��I�=j�S��y�� ή��6����l���ׄ]�I��xT_�S7r�QW��O����Tc���ۘ�b{|�iAH��A�;{�i#3�lG& ;!�v�'��N�R�7Б��y�H��7�����2Ւ�HJy|���1���ٙ�kG$�a�F���}�n�<>�T�Ms4�1^�SB���^��9b�5�S��7��x	Qg71��I�{���mGxC�1Ҁ���R�U�{��)W4h���<;+�d<u�&�oY����9�N�R>��+�^k�~B_�SX����ɞ��)0#����j�#� Sٌ���l2#08���ը��s��_"�H^Å˙>:�Ѻ�#�9�m�S*��4�֮��p�팏���_�PQ�܉�b��4�[�0y����ڜ��eT&�[k[�"���ߑ����L#;��h��`�A�F�+Œ��=
Eޑ�������#��q���vZ�i����R�q��+�f�����-h?��]�ja�W��!�%��&��e�	OXY����W��a6��"~S �S�S<�XI�&���cV�K,��-|Pt��%��l�n*nP�%�V��6�D�s������f�E�EA����~�����*lr*t-�v��؎7[:+<D��MGk�s=�kS��|�$���f������gH��Ao$#g��
��}_�#��5P�}���? j��Z�K�Mϔ%dDt��k,$���5��^�sI򫫑5{n`Fet��c�p��?B���/2��ؠ�d��x%����>Q��� �L���hC�A﫠���λ���޸��gС>5I���h����|fm���j�˻KZ�GiÔ��;Q7���hG�rf!�����ۛ��%:�_9ˑ��q�@��=��GQ=M  ��ˋ��b ߊ�8�����tz���~��w6��\i6���1]���{u�AͣB\��3%��G�y'��%�K����Ӑ����e�N0�Ց���e���eZ��xK��1e��w��ժ�9�ơ�W@ʢ��6�A[
4��N��'�2����dLp	�5gE�(�[Χ'��Ў;�+m"��P1A�x�{������6��X�h�,n<�A��gǶnFu�:%��X�� ue��o�6E�I�x�nnG����C��ir�(ޱ��]>�H�BC1���`o�Uq�S�8��n�*BD
���&VE	ةs�Z)di�`��j.5C��כpU�Γ���#
����7%[�������뫊@3P+@��vB芋��7��(�����ȹ�r��H�W}�u�Ж��X����8�e�MV��\��mm�!%_e#��k9q�(%�@�&�e%�Z!�86�5�U�;��z:�����}�sC�mx�hh�=�������!+�SnA����O� ^)
d���AoX�F-}D,���>��9v���4������z'Ƃ�'K=N��ms�K���t���0�+�no�d���u����%�@�Ũyn�/?K+��_���`�[����&�A;��%Rm`% ��ѼD��u�]��z�%�9�H�<Jn]C��e�Q�S��$����@,�S�q���R�$X��U�e"�w̮���1T��`2�EA�UB��$�7q�㸾�$Ҋ#P76ؖ��m�!�Ju�͸%�P*Ӆ0�:O�y����z�[���,6{��j}�q*�.s�Ԁ�L$��IP��n��8�D,U���
H�0%hH[&��T
��`��ٚ` �.ZD��K�ΰ��Y(��^��lo=�NI�u�Y�=�Fp���y�#��ǅ�����b�]��;�?ct��y�j�cN��f"j
�Tu����(��pTZ�p��+Xι��O>t�d�i�kV�C�ts��ߧ�:_�ͧ�2�0�;���5fo�k��������ٿ�X��}g���S�Tψ+�iM�W����?w�p��Y����\��1�;�K�+�����'*����k�b��E'L�ue��7v�
#�r�g�3�k
]M��g��G^���z��O���Q�\�h�áG�T�)�����a��uY?�ݼRm��7�5��8>9�?��:�$��?�K�.eGqt��G2��8�}��,t�{��W[���$�b�Ym�<���O�+G�?�̞�2ɿ[z���Z����/x��匡�4�a�]����K����7;Ì�Z�	.�A1_�?����B|�*m���#�K�'��q��>�w1��GFu�I>����01�j4ؙ�[b�&�D�-�d�g�w�A/���5#�	�/�&D�~�gPUn�߅/m*i'@�c�ӚB?�׮9�h�`Q3e�O�v�b��>n��t����(K=�R��T�e�ڞ�|"W�#- NG6��V��[�u��^>���f����q��\�UNiϹ^�:��S��6�M�qD.�6�*(�O���l�x	[�W^]�*hxn.������mʐ彴{� na��8�!?ٸ���jh�\p.@NT�
�'�h�9O��F�4o���m듊c����Tƶ��Kz:�Sjh: 'ÏL:���>3Ƃ���N��r���"��*݌���TKqD�o���"�����8��%������h���Be���6��_�ˋϣj�&�
�v��j#G�sb,J�D�*߼crz�F��q����F��z�܉�[��5��0F3�`��F�Mk�:��r���E�h!���*jzӎߞ�<��.� �;����/p�J���+mؗ瘡�)S��-:&��#=1/t4�t2]JGq�h�sO�f3���L{�v#GM��4C�Y��Z��k ��0��Jʪ}V<
M��.�d�FC�aV%QK�P���R��k�t<D��ݩN�X��DW]�7�Χ�W�B׀��%b����J���;�����4�M�Yf'�l=�E�G@��첀P���n��K��Ј��-���BD��ġ�ҽd	n�۫C���?�B� ve��	\	,O���������s�����XiG�gJ2������\��ߞ�Z=�N��¾�3 �\�+(�.�p���d�P����S���s��� �Kc{$\���}�y�1�/%8�������G���P"LZjd��[^B0��'�?43���#I�,*���&"�����Rå48Uʡ�F3�h|�� �#��/�t�ع9��w^��{@��+�=���e��Ο\����3��`��dp9�{?���7�T���8�r�L&gj�'�C�î�t��Y�t*������@W\�Z�Y2;+�Y�zd�4���Ɍ������W���5��Ԅ���֐�Eė[�s+��ӛ�%�ⵛ���{��Ml�u`c���p2q�F��_7��Ш7�rz�쏞��X\،Z�J伿��h��E9e�w{�Z�V���Hp�<�����^&q��q9~S�_�5�����ǻ<>���v�Qߊ�֞i�Ʊ3N�4��8,����kk ~���j򿪽;s�iݣIكK�I���1� ����v	�����2ˑ��3���vM�FC�$��7e�S��"��Nh�V�I$Jl����p5�)�����!C���x��6��z���/$����@O ��c>E�1pM�N��! *�ǘ� .��~��4����^��2��F�}c�$������BP�p����Ȝ�ց��,z�e�.�V1����uZ���>����;���}Z�̩��Ѐ�2!�� �#����3��a�D���,e2 �\A�ZXC��#�q�M���� ]D�����K���"u���h��P �S(&.9U��N8���'��>G�g]�h�u��QѬ��L�:W��?�w�oBH�dMUۋ�"�`D�1Z�T���#��+��۷\�D���3O���YR]-�;���S��Mk����6Tϳ��[����b:���2�z���!Д[w.���&x�O�1p��7��)�U���;���+�>V�Ex�=�9��&�ҳ��L���K�Uy��RO��-o�0-�L{��f�q�ln�6���,i(B����=>��À<�h��d$��{��Z�h�VR�f,�=��ͳs]��)3 EM��6�wᵝ��UȺf�έ�.�ji��H�}�
M"���ET�t����L>�>�y� h�)N���nט"a�Z�}ǒ5"/�N-�_M��V�6���Oȭ��h3S�qA�-T���Z��j�f�2X�i�t,��R���$г��ӯ�[3�M�fn� �N��ӷ�ׯ�^ڼdJdR0?է�[�ֳ���:�W���J��0p!X�?r�ew)zLWVF����$��o�}�u�UyA}'�@p���C�o�	)��!4��°�����T
{J�q$z�y���7h�_��J�5�~��*�P;wd"��J��U�����q�H�ned�������*�%=��!/Gj��o��������&��dh&��^�u��f;$����>@�� �G��akJ���@�x�.��������qJ~����4�6jl�z����Kc'Q��P�m=)�o�68�
C�p�v�P4I��^[&��ih������eﯼ�)WA�� ;]YWV��ٽP9Ԣa���
]9R���OMO	��((��3�Ex)��`41Pñ}:���=�,O�zhǣ�m�~�|6m��f��U8��tI�$�_c�hAxFC�&Q�L���^�����h�c~����� �s���N������q�ů�7�u���.�%��xv(St��X
��=i��?�����Ց_��1���MPf;�q�qB=���,{�����cݢ�9�Ow�&^R�`�sy��~c�詃�$�p�p�픀Q��(��ʤA���}-k��r0Z�����[����g&#�ٕ�n�,]�#�xeX�5��jI��U���\��\�`���m����=b>�Y��Th���gvX���0O���hulp�y@��(�{JPڞ�bU�>�.�{����� ί>d��y��"�������B���"*!�|B]+�F��K���&!�u��H֯�q�(�V�s.N+�q�O�J���������7�����\=R��n��ݷ颠�����
�:8�I��s�ż(�L ��xM!PE���Sw��|@U�v?Ӯ{��XTe3�7��ܪg��	�KE����ou����(�*&�+"$T	��>����W�k�Mw���ȹc
*���c�	�L�%��_����
A����߃�V~�]oz��[�J"wR��>v���eMN1Ϊ�q}�����Bƨ^v)�P�^x�ZO]�
��~N1B��Nf�h8@�@����X�ڸ�R��B>t��9�KN @䟑
wMۄk����<jC��pX�'B�0s�A.����_��2K��y�#=1��g����������ud����#�B:�������=����ۖ���8���>��(�[�!3�G_pl#Ҿ�E)[��m&ͅ�ӬYR͵��	�؊�c��i.�˛A�|I��C�W<~c���j�|z���مC+Y���5Y����i���ԫ��t�l4::/�an&p_L��pq'����up�<��.ߔ�Ƅ�]P��1c�)��fO�n�g���`�E�PG�Zm�1-~0N����2�WYCPǻċ�\������ dG\�/Kk|m���XǺ��@g�iӕ�UxL���Z�h���ME��H�iA�q� 3m�ٛ���pϓ9�O�|J#�r����PĶ�3i��p߰\,�z累��p~��F�&i�GS��"x�&�#n")�JK"��Q�nF�ҫ0v���7�:��f���^8��v�2�[�SC)���h��
��6�ҡ�\�.g��|n��h���V��"�#��0���,D7𝆦�ZA��8���>8˱0�e�h�ut�]���J�ұ�X6-�I5p�>&Q���^���D��H�B$������:u�eeNѪ�b�A�|p59��،?J���ڢ4`��OU!��楽n��%H���7n+�p��|k��ѽ][�����y�B��({z�ڻ���_�p��*���F�c��1��ѻ����	߽�J���kC� ���؋����՜ח�o�c�p�V;���т�����*N����-��M������lsO��*4�B4g���7�bY����ܖ��Q���b�����E�c�v6\����ih-��bZ�]e݌[��Sh�t
��aP�������%�B����B%b������T5K��co�Qu�e���,Zm��|0i���/=z���MO����F�,�c[���l56�g�_���v-�
���0�4�]ә;k��y���R�-�w:r��y�%!�"�ϐ(d=)�+����H�蚚����ޯ���ˌJ�ˬo����)UC���?��n ���
)�����uO�}}[��~/���Z�.<��
�J��캃4ht�ݖ�6�Ed0_۱/g૩��c�>8Q��+���������Fk�$�|ǳ�#�}���1u���� ��5(�a1��	2c�g�O�"j��M93/�*>�C��j>���{�O^�I+��I�L,3��T��E�*�E��"�K��ԇ���A�����'�Tk°��fkVdB�>E�؂�v�W�^΁'/�F��q�K�m�lf�p���D~����W��W�z��U�����;z�V�iIv[����t�����q���*oڶR�E�P��b<Jzg�P������M��ܹ��֎W������	�# �_ ��ҭF�J��D���+~V������ʑX�!u_V�y�5��nP���h�NCfZ#@�Y��K3h� ����
��k��(�ď1�?]�����l�9�9�n�V���527�+ŀ��ƃQq���1�TI���0ԓ�#���j��t�?�:a�������}�Zj�^
�M�)��T��&%��:�Z#��>L����h���[0�sr/�Ih���¢��|���x׆��3>x`�Z���~����(+S�6D��5���:Cv"L��NPT���3PN^�h��1�j��֣
Y���.�y���o�r��s�a�o|W���O*�O�;u��x+���4h��dW�5�E8�m��5q���͑<C[��6���'e�D'SV��ѵGS����e�,(��(�Pg�51
1����k�rY��Cv)�������ۺY��H_%��r�>�ZO��0���L�v����:b���>�6z��7�(���g�˓�U�e�E��Q�{7ߣ��B!� ���LY�!EK�_��X�bD/7���.�{3�/9�m6�V��'��u8<W�*6L� _��,τ��I٫0|���4�0�i��!,�<�9x�B ����H�ܦ�\�D>|��qk�pa��Wj���=�ȭ�]=3�X���:����P��P�?�EιH���1vnc o����M�t�;|n�}���ƱtV�Ԯ��hF��PB��P>�6�����4�G2eX�f�֞{�#0U�{a���W:5�+,Nj�هΗw����࠶��YuaۓZ�.P?р�1�0�����7�K�U�V�_ַS�����AV͟�Y�p�`Cȡ��2��JҌԿ5�s�X�ͪ���*�?�T�mmt�	8Bt��hS9��3}1��Ij�ݣk�G�f4,�%��dm�k�KH�q7b��}��AX�e,>Fp;�.����&���G�8�s�%O>����&�����:�n7�vT`2�sBX����4���/�e�U_��$�/=��H�$~Xq�����7��aǇhǍ�(˖�ܗg��t��!�<���_R"�zg)�j���t����F W�0!hק-�ǣ�@.�;	n�2\
�x)�S�iĿ����f?I[��\��%�%\�R����^��-�Ce�A��h�����7_�)��0ǜ��R���\�F~��X���偰��V�0_A`��֨�;��N��jkep*���%��P���vRԟt:�VI���� ��>l�ŋ@/�0��4�������U�q��1`I�ٹ�-jQ9t������t�BD�5,d0���DF�u"�CRJ��f����^��V-P�!wJ�aL�����+���	+5ޮ{���n��4;�dujF�G<�
~�iC8��͊q���$�)�T�T�JM�����7V��hk�/��T'���1�6R��	��{s�V����{*��7)uN��R���{�L�T:� �C���aL%�b��o��!��d�:�^���X|���ɬ�r�`�3��Mi�U���V����4�{��8��0V�uZ�a��,pw��S�J�O�|��F�<S�:�eOu̾�~��iVgH
�jRch-���"�=2���X ��y�(�ЮVZ�DI�b�2�M[�hOg.j�eP%o2H�)6k�m��sy�7�N�T���ν�q��׽�5�H]���5@���w��jO����lzH|I?���Ȭz ���Y2@>�}vA� yaγJ��q��g�6%�`x{:�`��Xz��.�=�
�ޠ68����\��2�U��J8�ta!g�t� ,�=e����)��5I$�3��� ๎�5����G���	��e>�p��ĶQ�pL�Za�Z��ܢ�=��G���BPXO��<�ć�ÃNB!4Z��K��Z�@�������V��wa���eo�n��X(h9|�.�)��Pw�{���{���.Ry&�X7������+�e���5��𼃕ނ��y�׵� ҈f ~���M��h���w����di��+��pI�-,K!�e~��g���v���A�6����y�?햻��C��\¶9�".�E��R uX�aS2),�5��p+���y�+-���M�=��׼���wG�`���5/2�J�k�l�z@V=PӮvI�(?���v�����Xu�����2'��3���]�IU8���(Gt�߲&;��wͣ�r{�b2�����j$�}l��(�
R��M�jd0���Ѵ3�e>��[w�M�7)*�q|�j:Ŋ�������v�Jl<s�32Oa;��-?�uUF�%�7ا�~P�o��������#s�Ȉ30ʫ��v��z�Qd���{a�Dx��N�#Cw�X�_*g^��2$L�����j�*���C����}�	�&g�K�*zVC�j�����r�̭"ɲ�ѱ.�r��k���#�C�y��."ձU����w��!�����2=��n�d:H���-��3�1 � ��_yLY4!8�D�P�V��7�#���ᆦpp���+҇�E&ک�2H��<Bj�-����=�3�8�LD4?�'�:ߘ�^�È�w ��E��9�����n�m�&~���p
r,/��:R"@BW/$��>U�XE�o��܀#���F�t��Mc� ���D4�ƙ�mԻ؂�Ie���U�Sz{މ�_�8�t�����5}#:`C��9�'M,j���K*���;\B[0�]|��>�H�W����.��ȒV�A�#q��{�$�T@W�rʖŕ�_zG���-���
���.�������a�݀p��m:m�(A7�d>�	���x��]������YD�<���h�PH�D����Λ�L�{����F���C�K�֛nV� ��j�͜Y&2�d����HDm�n�0��4�
��9ц��`}�ԥ��U��P*v$�s6�g2��TD���K����Bj2��e���3��Q�r��N$�?���CM�l	{Ʋ	OF "v����ܜB����H{��X�������`!�vEv���h]ׁ���^Us|��GN�#`|I&+x�)�~�lU"�$K�P`�4I��9a*�/n1��c=eZ=Is2�2wxڲSf?�l��6	�S��Y�3�2�G��0�H�0�?����.����H+�.����:��vZ��@�K��Vxo>$ď��� ��n�x*�(t� %)^qi�:��7F�g�y(/Y��#[�'x1��5����2R�9 � ��[K 9�am��1֡���4Z!	;�
���BY�������RM���v�A�K�q!_p���|�0�S6�T��0��`��TN�i�鹵�}���%�.���@�)��;��~��	�h6�}G�nr������YG�����qБB߯�'�/���$Q �E��(���.8X��>���Uoov�i��r���v���.��`�kPh~5�;i��F�m��y��CI/⦮��|/t�\,���[�N�Ef�xWv���Z�_#�g��D��1qq�Ǎ�nw
1t�Ew�f�[`�½�Xg�wA僑V�x�n���и�*5��Ɂ�cnD���O��+U�pO�:�ѹ�Xw����%w��@ö�jl�rC&*I	��u뛫��]0G��G�̩޺T���K��/�����W�|J}h8b�CI�{���*��`*m�#DW|��H��Q�˨/0�I���{g�&MFktV�m66�_{v��`�F"�T��=�Qc��]ַKy���l���]�ʿ�0�E|��+�����b�["0`���*��::Emz���M��~]4b8�Vy�	��M�7�b�-�0�Ă����K��7�ׯ�|a��2�z$�^D}�Ns�&JL�v;nvD�J�1�\;����^u��N�I{C��*����+��kY��v�X:�
֎��rT1�n��73��{s,���l�^cA�W���9�3W�i�.���`�������.Sd5a�Gy��ȓ��z�(�x�C7�i�b�VE/q@�z������
ZXi�43�8Q��v��Ұ��R��%0�%T4�:~!埙����鰺�cȢ�։<��䓎(M�M��C�Q�NgԈ�J
��`췫�̙&�fR�p�l����B&��Mm���D�_�dc�3����$�o���ҋoX}	n;=�t�r6 ��ͥ6��	��<��h�%0�ϣ/BaM��q��#\�W�9�6M�t��E��o��r�,rF�cCp�5�w�aM=�
�-�t�xU7T�t݋��W��$'�ףRcvR�a�P���	!S*��_�#���F��� .�uyM%��e���n��7��B�X-�&g(N�a.$����u(�;/��cˏ�DT��.�P���a;�Ҍ�o���Xȧ�S>�")w�w����%��>�ا؉E/��d#4,�M_�fnN~��@�ْ|��m�-:s����`�,{h��Tj�<#�;��SDY�#��j�����HD�vq�l�G�CeUCCd!�e��l���~-�3��^-'��0G�x�ۄO����6��_Є{���}���W5�%�2����nq.�94\!p>���B��'�L.�@�����%�Ɂ�	
Fn�w����0���ED���<9��5k	m��+�6�_&:%�͗�A�ɂq��Xc�Aӝ��!���?=�5�7�I�?� ��Z��2���,&4�X��]8����G�ȧ,�/۫�IB����
���[�GGx�X^_��.51bw>���X�`��R+N�U�w�1�ޭ�ћxVC�H�L�*�+��ȭҾ��dM0��<���!�-�	\�bL��F�"�%d�$�ю.��^O�Ox��hP��@��|�C3QI�ow�g��˭WC��8|R�����U8��K���ʫ�����ມ�W�s+@�!`�������C�gE���Z�#��nD�����x�W����z0�>C ]�J�˓�Q�	+�R:��7뉭�A��
`�R�Y�H�d�s+})�hՙ��'�~E�2|hs�q�o�!����ܻ`���іgL-�t�GA�k,�_�(�~�f2#���/0]�?@� �&U��;�7TN���j��N1,�S��V4�/���b}�z&_s4��9�.���0����w0��Ǒ∟�Hq�q��_t�7w�
���%��x稆��p�#�H^�W"9�3�n2i�ڛ�/����V�K�l/�݁�̈�(��p�G�­�A��&���B�)f��D��в�N.������n�WL<P5*�10��r6��MID���u��c�|�R���65m�`X;!>�DU��E�\k��V�6#5�P��d�IMy�Qe�e�o`
��8��	%LF�����L�JGZ��)K~]���.Gq�*ه\�����L4EǪ���/�O���
/�����!�6�n�S&S�h����ca�{����O����"��_ t]�򰶜I�I�,� �a?���;<�E������w_i��)�[����^^)<gVy�J22<|z�J���rzz92�ۣ05���R�X���Q���y��-��7�Ec��2�U\�i��*�Z�!8����k:�ٸ��:��ᒦ�bx�`ڄ�!�ԁ�ȑ(b�fШ����9!�ӊw�7�7��6! Zlwp�(���4~�3&����M-��K��zI�/���d��K������H6d�4���ĺ�u�k:�b�����{���O�T�-��$ ��)�b���@r�^|�"/<{md�|�����W��:� ��Rf7�H[oS��9�b2.���,XK�`��-���"8�Q2#7�{w��ن�X[�X���z�;W���p>�>K�k	�*����
��.w9�����z��Ub,.i�S�.�ӽj���n����Ke7J����c�P4�l�t�a'�|}�5���5�I�M���*��q��iX��F^� �:\�"3��M\e��.xjֵU���s��q.���b�иn���?!�a10��<=�6�JTI�	b�r?���w6'���B���憰����k��f�"4(L�R��US���؂�J��w��V��W��������ҵ�j�NXl~���2�ȡ��U(�+�rזV�d�.�ƚ܂�"�4t���1�P��I.���%s#��0��f���(t^��nbT$3�KM��g	�,Wطޏ��P@�Q.W#u��cM�~��p��J;���R,���Y�'���h#E; S�ǆ9���,����I���������mg'/��w��k���ٿ^�E��^���n�l��_��F!���ֆp��,N\MJ����o�"a�F��7tT=����	�$����5~g�j�f���|��n%��1P�\��6mQ�dOk:�%����qM/#L�3���e�}Lc�c�c?*��2@��s�.v�0�VO)?�u7���\A���
P���{�l�ą���'�hi���YEgV���0|j��9Y���crX|�x��ԑ�):r�U��r+�C���i�'���8��tPu`١��ҍ �	���-n2�A|���ō�'}l�"�y��߀�V�������[�@�g *�����$�t{�B��UD������V�~e9s��b8��d'��YH�^{J����9�Hw�'
�8�d�,���:����nj����/��ʳce4�����ܞ-�k�4���U�0-i�Y��Š�Tn�TS�t.s;����qfK�d4��<�U��6kQ��7�eL���0��Y
�������8DVZ��]�������c-��8�Z��:�j'�t<������ʎ�S�?h�|nMע�%���i���M�?S�n��E��۬+L"�-E�W{��m_�%�Ia�9;�E��5>%kF�w�ՖC����UAo|;6�%�����e��LC�k��y'b:�	��r�`~1Y��\���k/2J����c����9V������
dct�߼7��RB�.�II���D�ŰcҥB���pڂ0R7�V��Y�@t\�/�n�J+�<��j�Rr�̩�����6�w���������F��$� q�j�F᧸O܋��E�7�Kg�܇U"�C�1)��P��߯[x�!���;>��{��Lw���&t��l>X?�yl�o?
��8�d�!��C�8�q.e1�vGcY���#	��e<P+�}M-�����8?;�`;�$�ӣ��C�Q��^W֐�Fn�]Ѽ������ϗ6$���;ݐ�ha0����o ��Ȼ��*e��ר�v���`kgw?� y�<5���I�J[�w���ϊ
��K`/w���� /�,1w��=��I�<5=�tEM�W=�'��	>&�����>�慡c�k����m�.]�]���u��FyCr�3��b�u��Ԓ�պ�r��ԈgR���)���R�Duا�F�R&#��Q,�"���f�){�l�5mP��^æ,�^��̍�LrRI;��bq�	~��Ǳ��N��)x�xc��Əd�iZ�T~�>&�n8(�z��HO���r����~�r��J��쾏��X��
M����Я����<���f-����$��Z�[A U|��Bf�1�б]��	�RլT#Em�����ԒB��nz�l!	I���;?yY��q���Ԁ[�Z֋�BF��kGo��"�A�ּ�F-g&g���w|���m7x)�R��3)g��F|��u��O�(�r�������M�M�H��R@rMf��Ojs3@��L�.?��)�f5�~�OO�#�=
����}��H6;P���J���? 6��8��U��Hݦ*�qM4,��ZѲp��1��nQ��_w�b��ظ��_͜/�Ndmc|�{�<aw�)!����6�P���X���|E{���E��\�
�%z���5��.Q_������MsUk
��?:~��;KR�[vI�e�F~��F/�����X�6��P�;
F�K6�B���2�����Q����D���w��T�X�-�1\��{Mtq���X�9��a^{X�V���F��`��	��'y�z귅#C��Yo��<�Z ښ&�ek&��|pɥ8�������_�+��|1L	���
�����Q76+���/�C�U[��NZ���5���3��/��P�U?�"c"��
��<�|k�Q��s��X-�>�k;�o�|�1^�)���Δ�A�4�S�"��j]�ϩyshc��H��g��R�r�)����z�ۜY� D0d�³�r�/�rȱ2�+RX8����g�/��v�&��D�4������@���x�p/�=�:�xi_�Ѿ�Wy"��[�ث^W�c���iL�`���@B��~��-?C
g�q�@�E�	�f�I�ո���x��#��4����C�ȟ#����	m�����0�?�Z
^ ˆQE4�&�b�!���=����.��Vү d���J,�;39t�o�.�
+VD�]��cד��dH��#o!{)|@-���"��o��T��D{�^�Q%�%���\�iE��	�#eUàWZ�Y$O�5
Hn���j\����Յ"�e}�s궟 �C��&,8qy%E�3%;j8�*MQ�)���y��>������ZAR)�G�"P�~��	Z1%�p��Y��< (���3QҢm�Cu�Ong�@�t�H`O깳��=���3���T�@"�9�<�ƾ��ɭSv8p�pjZ9+�{|���"���h����;#$ͷ4z���=��Mp"�;א�/�ґ��$�w�]�p����o���\:I;k������>�G�xNT���6�W��M �n)�DZ-�,����tgr�0�,�ޚ5�D�ۄ���-��0b�B��E�u��
�=w�*���}P�p����s���_�����_������gr��<��xrX��5\d��8�WB������nZ�\��h�*� |$�`V,2�sʕ�̴lO�ҟ����>Uh�Ms�\��vN��ݎ#ft����C�H�*�u���Z+2�*�|+��v�+��f�E�M?v�b� ��x��z����p;趙Y΁�;���9}��Τ�s���]��',��dJm4�(��b�XM�ۋy��hv���ӱg�L��+���C����s����VGM�V�ɱ����.1����A�C������~�`aD�uŔ�b�ȑ\B�����5A�|���L�V��&��Z��"i�kM�}�eId* 3��fXi�0X&�'���O�j*��b�栢F8��(�q��#��O}:�
��mI�C�L٤�f����Q�� ~xa�o������T��&0�֮��`�6ꀹj$��l�)!4o1F��x'|MC�Kl-�[�k���y�_�5P8�l��2'�D�q�׀,
nBZ @6�k���~G�N)0���
�-S�F�����R����ĩ
)0p%����v :k?U��,�k��z�lYw�V1R��-m�C�Q�O�:aGws�|U��*�1��Gi���UA�xe�x��L��1r�d�3*%ԫ����NK�y	����F�/��]j��ݓ���I kh&�@^�����Pw��T�Φ1Ō�����*&����a��B�E��ET�|�ғ��aO��5��6T�P���3H1ҕ�Ϫ�΢<���`������H���a��@��q�2���������|���ゾ�sK<�҅6�K�♈�9����eG�l\{v�lC�3��w%s��-R\��:�k#��R9DH�C7F���e n�����Ae�Uh�����E4Z��o`6��΁��jՅX��Ul	YY�̊�'�io����L���?;�h�t��vꎧ�n���-o��!��bL�w�Ե����62�9!��!Eݰ�y6�4� �y����2���U��[t8�ř�Ŏڻ_�Zp�Ex�B�ݲCi�s,~�:Cx�(ic�g�ק�Y�W@*��:4�s_t���t��\�X���w�A�}#jVp�5��s ����zސ�Ǽ(����<�q����y^X���B4�AO bQQ6â��_�`���潶3�
=",�g�򄓑���v�/xMR��k�'!٤*�r|���u����P��6
΁��`�g�錖��KHH�R����}qt���'�q�N��ra6���`v�����w��$���J`��u��U�Z�=�4���ݜ�Ͱ��>��2n�^:�����;��u錌8��p���P�&�Ï�a�4��m�9�k"�r���20w�I'���wЫav�oӗk�7�uoD֠�M"ϼMg�wD}B��;�������8���Hn�$OfuĖ__�Gm#6�3�[S��R�o���+� g������m��7�j�N,�0BuӉu洉�T�P�fz�'��)x7����*�o����k�\����%k��>ΐ
0cp��zRQW����I�L Y��$��6���θ�r��1f9Y�.�/7H�w�==��M�)%$Z@;�@�2�<�f;H:_���+�g���GC�l��H ��|dVpEkٜ�nN3Tbc�a��'�XL��"��=���O7�L0���q�'ԋ.��/Ő�ԣYdR�Jѕ�pTH,5������"��-�����ǳ��U�J�|�9"�آ�3����@;�[��h��s+-4��e�mFlʔ��*~���ZT4}��P��S�C��M+Գ7}*D&��.�1�6�:��ZI�-�Lg���ŏ�h��UΖ$�ƶs0l�s#�����]���ݘ�1֬\��;Z�>�t̎1�����~��=���Kx.�l�A�2��4��I�kn��>�*XQ�U �[W���E�j�S�'�J��JR���'=��Y��F��P�8��lV�d��L[��?�C*��j�)'�)��Z���J�Bd�ِ#�� ���%Ix	�Q��t3�{Ţay<�e|��'��u�*�����eeH�(ךE!�s.��P���A�X�T���'�}@qÈ���"C�z��?��=�}���i�|�k�y��<�/�{�a�G�=��bz���jw:���29�kGK ���9�� ĸ�W�y��8��D�z�G} ��6����T%�������k�����+����d�Pa���f��ٮ,x'p�s���t[���;��t'��C[r�Ƨ|��\��R-\'Ѿ�5�b��eI[+�@B�̑NUx�I�&E3�Gl����7��	���	��nG�:�]Yc�\IlX�{�x�3�l��`��Z�^����D�����.G���"��d�~k�����R!H:�؋�
~)������"�7����l�y����[q�T��A2e/W�N/��ث^e.t����27�{y���"+��3Wg��a�x���#�I�V��(l�8��$����6G�t���G�0e�)&#q�\o_����
A^��xK�`��y��-��5z�n�~Ɏ��c��8ʶ��f�vU��'K=�W����K���>�O�5�&�o�-�K��O��4HBԸ��t�@���ޫ��O��R_�ڙ��|�PF#���5 �l��-ƺ�����������9��?��o��<q�����U�����m�k��MmQ�'�1�М��n��k�� ���mn(IҀ��8W3�bĤE*��ݺcal��F�T�jj?Yc������_�b�en6��W�jL�|=և7��AcgS��ͽr��d��D;�zĦsKzF� (�sr���ä�* ��Lyw�*���.�m�䅯¦�#m����;<�����/�º�\��w+�Ga̞B9�T%��%��P�_��1Jk=U�"�5���Jt��i҅¸zb�c�zF��-֔S�T�(q5�Xĵ�]��^��/�Xp2�a~���mdU��;s���nS+^���)�E�ВE�1=��$�=�!>�Kw&�R�ʷ�싉S�?�B1���zR|
����\�O|Q�Al[����k����c�6�4yR�f���SN��h���v�8l��=�xk�乒�ƈ��K���z��4~J�޺���(�s�|}^"0����xYڝ��8�&���0��� �. �jA��#M3V��.�x�N&p{��\(jw�ڨD����5%f����� �_+T5!� \���`�J� H�ir��Z��ļ�8�����I��|ՉK��x5`{����_]��}w[��oz�j�݅��5�r��s���K��ȅ�b�4�!BEx��g:�ig��+�	�%�4X�6Gz;��!1ìY���X�Q)�WR+\CX�h��{���k��E�`-�D<�8@�V8>mػm���=�L7����Ź[�2��IK�X�KA�4VJ�U�E��h�He�P�U�X����l�{�����h1�cS#����g�ߙ8*�PȱQ������}�i-�r*��㒣5�#���2��2W:!�BF���$��Ci�j������C$�)J2=�SN��KNsm������=���\�2�]��KK��	�)8�>(���>f1�055��J�E�E���P��y"���"�m��[��[[p�ڨ�k�=�ʠ�`��"W�� �/饝|�Ý�&�Q$��]@�r�ӥl����kD:���8����S!��w�o>s����äG_+�gb�Ծ�L#6�pL��^��zD =��U��_��`~ݙr3�|���*e��"��m��}0�k˂�.�cx悋��B�a����|[Ht� W�q��&��X�76d�s͘e��rTQ`D��M�<�Q<�0�[�yX��>x՛���Cj��a�%:� J"����PO ƥCp�J��4��M���Y�{�pK�y��-D����/�{��*���o�r-&��14�H%n�ǩɰ	���|l����z��X���bڅ����bF�R��b��^[Q�����5�f|�Hy(��X\��|J�,��l>�*�d�A��υ��r,in�A����K���tG��������3Gm�
��+ʙ'��W�=�r�����ɉp+~�I�!W��� N�1N��0��'Z���(jdLA����	`DA����P���c��Ċ)�+���0�`#�R{��!��G�9Ӣ�`��S�6�(�ϛ��п�ʟ3�[�	�lc�N��~-u���M �_@b�V�F�z7����w�a㣙�F���r嬎��/������*�Wj@�a�?`88�ʜ�A�qǄQ���rgF��sFW��j;ۼ�/��)�7�>3��
+( NoϙB�w:��`���ݒ�|�R�2�uq�-7�(B�Y*�\KUH:�(�I�9�兌c����5������nu)�^8�i%-d�v�/F���@��׊�2Ȥ:��Q����ȼ��l��m|R^�b����y����6�g���=I�0ų�>���n�~`�#��e�_c��ل|k�ӽ�3�!н�2Q��a"���I\1z��6al�T��)�a��Y3��X@gp������4Ú�l�rN+��8|�)�����M� @)�����|zs����=��$z���-�s�� ��*'�Հ*6�e�݀�h'�RtR3���=�ޫ�����37[T�,��r<�p�`���σ�Յ�Q׷�-6�xR-��.�=� �w��	/�p��ۏ����&��V�nH˽D�̅J%��-�����"�:p������F�v<}*�ȇ���s��zsa�Q�1,��;�1o�lbl<�Lnj
�ӻo�æ��%ݳ�'
E�Ӌo0j�cïx�� A��*�G���DƇ��"T�.ąQ�&�����y��~�cm��!���
��c��qJ~��`����vm��o�O,���R�h��oFS:�Ņ8n̫I~�#�FC׶����$ڴ��&�F��.�,��IT.������PqO/?�ٜ�6np��\�ѽM�wn�aB�K���NU��S���������~�"��9����r���Ĝ��sH����`��BB��xAg'\Ì�� �>�1Eߍ]���fa����>�͇��X �1�~�DU��mXl0��$cP���� 4P���QP�r�\����8�jo��oiv챒ڲ[}����^@�s+yY[:a�Ac�q�@��m.����e�uO�`�5�����7x�n+��O8 ��&0��R&�Bȴ���[�jLnZo�q��\Fh�
�7��&�ms.fzm��9Y��~hg�T�|$%��qA5�d�D@9g��Wh�	�i��%ҝ�9�� X�����֥.!T�^�\j�>��[e^�����3U��rb��"����:���B�)X���|S']�GNw��Kߞ��t'q4Lnl� �|�����C�q�m�n��_�zU��qb�_�ó�J�F�"�8b�SƘ���bd�5#@���Y�L��ÜO��wU��l/\q���fac����3 ��b<S��������	�*^��H^������Jܞ,���_0ܫ2�������2��z��+*U��/�K���d��-� ��qU���`�I.�Σ(��&K��E
Ĩ�\ޅ��k}!#Ei�ZA������7���X�Pk-���;�/��A
'���ݖ\�D���%�D�W���t��XRX��λ$�G��nS�`Q3y"�,~�@�PW<9�1u�稧*�^�_�_(JZ}H�R�A e�!�@�h�x������9[5"�z#��d#�A��O��tR}�%�9�^�c~Z���+|琝�myq���pm*E�妤�z��%~o�������$2E���a#�-u4H�}�f��MJ�餿��ba͛�T��t��#��v�,��<02g�LA�g/Ӳ,�#LЌ�)�{R��
���h�l�V�7"x	�7J�y���p�>��k�hry��kнH0�)o��}��0t���#�F�6._�/�u{�H��D��p#�N�.�5"����r�HՖ^剓��ø�ߐ-���QjL'N���!���q��352�B<�j-G���j/��z��+m�n71 �dȏ-�rb��$��m�yAY�(��Q�u�0ض(�������p��{G�i��9�p��A����sdXu�J���*nYU9�0aOx5���i�a��Eۍ��ջWZ*G��U��y�2ؘ!�_���E�TՐ����-0�<��X?��ۜ�*}"z�#�I? ޲��4Q\/HE���K�ħ�,Di��������z�L_����+��������SP�ի����?[��*7spu���ucͮO,��S	aؒ�:g�������������<�:�4�|�a��LC2ʭ{Z�rm甚
}+L)�zT4����Nn�ڟNU� ��c٤�}v���A��W�v�g�{��0�pۆ�36���XZӚ�(�4r{Vo6�\c8�4�>	 }�
� ��[6��8D{�&���L?�Z�x�COD��莣�NH��4�9Y���(S��c��i���R��_5)���|�<�OOP���l$��ܸ4zx-�?Glb�����g�Q��|T6�9N\ E*0EW���d��xs#�1�+��FB��M�]z����}�sG�i�uB~�@4r�L�)ZI��P�0��j��>��z(�:���:$)����sxk�F�?gI�
[㡵��ͳ�gw��@=��T�9��B�' r���fug����N��o����n�����z�[�ͤ#��t��E1�sk񇁉���NC���@b�!����5�M5~;&®�c*�z���!~�"�*Q(bf���r��\�[�'�x0��k��E�,�`��O��Dz��(�K�0�I}=%�4��}~d]��@7�F`=���5pb@������!��� ��ŕ��|Wە�]q0�k���Ys���-ro��?����Ӯ�kv]եx�F�2�XY5G��@9�A��r�gr�F�	ot��u+��5_~Oll�U=�9�n����|�[8�-[��{&�|���D/aѕ�^T�Ҫ��I.j�*��AǓ�-*���	Q\Y �t�f�:�ˢ�<��S���;�ـIX�<]�pSi��d���ס˭�hF��y��e���{T8����;&�'�"�%ms�m=>��ծ�L��@'+y
͢B�Ls��zM�<<�<�Qb��s�'H��� �s�p,�B����b���J���֝�m�^j��Z�s=��U��yQ�V���h�.��v!G_�j����o5CIZR<o��#b\ 2bⴳX@ ��}?�Ty�����>���FE��� h�h��kޫ���k�Y� �8W�r$q{��5}Z�$��TG���&|nr+���A"Z��Qq\��S@�85�X2�F����ҫZPm��<L2�ek!�y��P���)�%�Y�*M�7jԈ$��[��v�E%�3�1z��l��a�0��T��̄b�7u��GT�̗��b1(�ٴ��5��J��%����g@a����HT@1;�*��b���q/�W�"����-*���d�n����lC\�6�ί�dPz�F��ci�.%L��Ck��	����Ȣ��o��
=Aƕ8�����8hB��6\��I�,�ԝO[752�J�������){f��bߴ��d��&1�P@ݗ-������G����*.җ��4���ђ�l��hP�Kܞaz�x��̶�p�v��uNC�.;��q3�l�y���4�+>-M$~��aK��,q�{Tb,P�w�!�{�����
Ҵ��a�(xg4ꅋ@�f���� KE��p9D��o��o����ځ�N�<�^��v?V���A*�kwY>2�O���6�M]����d�\zt;O��8�#�ǕJb� W����1u �`yd7���-7�h��]�9����8͞P���a�����F~�ri��u$�[WK]M�3#
d#�{pg�����i}�҆2@5�e �	�D�.�|��7v�w���H�'1�ϭ��P�F��"!��-�L��;|�gĦI����zp:�G�z=���gR}ϐ��z�_�0�俟(=w�@^��(8��,݀F�~�P��ém"������o���e������gS7���)8*�w��n�Ak�NQH�$H�uR�x�+��4J7!���'mHͽ+��w���O�}������Ĝt�S]:w��z�N�>�ƌ�~�iFgp�W5��WcQ�zn?�(���ҁ��(4��>�$���%��U<����g�j����Y�����U���n�x�4ݴ�y����H�.�J3��7o�Z����oę𬸃����q���Ml�!���#C;��u�D@��oFˡ�m�~EUr�M�)�MW����'����+d�jJ�o3I�����(��hҰ�8���]�f<�����
����c
l��������J<�"��s~���E�V+���έO<)�b��ka+�Ǿ�l"�"��2ĵ�uݍ�6�q'�V�0�:ь�/f��`�0#�蓎�	�:�8�>��*�7��n�����X�P>E�	�bb�j��Y�
Bgz`3�+ǚ�[H7XQһ�s	|~�*a�j^&��gR���]ԋ���� ��Ձ(ׇv��;�zW�Ư�W�:��)X���Z��$�U�RnU_.���6C��#���󛍈�i��LL/����F�f�fj�Q�A���]ZR���"e��m)�Ҫ35��QIE4a��jZ�}��пNT�4�*�tӼ�3�E)�8�BX�>��C�j�[��E���.�}|�6��,��"��L���n�o�׬/��q�G�X�ޠ�[vI|B�A#��,��F��a3��k0e�"��*��	79b�j�����b�շ�#A���Dk�l���Q���fP�C;N?�J0��<�=V뫻��uП�,i�\>�{x�B�>�:Y������0��yn�qޘ)��������S���9�e!s�:��]��m�����H�/�<�[KPA��%���*R�kh���s�f��%g����}�ӲWtb��2�(����������,@!iQ�(�%��m�8G��1���Rۈ��W��0� ��ΝM�A��a�jF�QlR?���)R�����:�o̡*�7�!W���u��,p9]LU���:@�K8iW@1�b�g��J�\[�	�{�d��3��d!��-����=�N�!���W��> �:<�1o�c����e��$h�\�D�g��-Q��A�n�J�.�Ƈ�����9%�4&i�J�m�䯆��B�ϨO8T��3�/;�!p�ξ�����̀�/[���U[P�*�:	�[��~��I�J����@7h��x�2B?%~6r4�X�+{R��Dk:f�9.p�I��:�;���2���dz"��仿�:h�p����h�e�Z��ݗ��3� U�'�>4�Wȣ).-,B����l׊}I�e�w�>A�B�A�KT˞���	�,���J�H,@I��^�HNU�%�}�1�>ԤEw �88�q��I�8�4I�����O�� ��_d�q-&.J��i���ɸj�,�X-�|CL�}ѵ�EilwH��,����:���B��A�HE�V�;�٘�7ٗJ�˙nYTzZ��;��F6�Q$zg6:OJ��b�Hx�Vu��$��^��?�y�$>b�TWJ������-�����4R�LO�v],0��[?��V&j�O_G��N3m҈7|�o��
SJ��i��-���WL��7��YC�e��|�=6�	�!����P����N��6�²h�Vp��Zl��kUm'`�:.�8TV�ð�7S��8`�����_)��E����>�s����5*�a�O�5��b��k�gi^���6���5�@f!���v�^s&�0��&�F�l�_����H��2�5�Jl.%N���ݛ�v���]p���w����΄zJi?�_����|L�s��f�N�:/��X����r2��d�(7 ��I��b�dN�M�h��L!aS�s�y�2
� ��־7i��j�/&����<.�;:��% �Jwr#�b��J��d'�s��J4����z|�QK�����P����n��.�B��Q�_"��y+~@�`�X��B�3�JZT��,�g��7�B�]�K��D
�d�]�]�鯾~E��J�@���o3���j%/���o�)�v��q� �Nj���Ϗ_7R�/6��(�����|���ʬ�A�Y��`��ک���g�gr�{��]B��ɛ�g�����e.�u1�eP��i��lс���2�{{�����&��S�S�[W%�����k��*�v%d���fO22�ܛ�:?��}$��Iv�����'�@�E%~q��,��ɵ��+��/���՘�ly�u�uh�y	�b nE���	����̧��������F�@����A�jk��;�`P�X ���M7*o��J�?T�)G�@w��p�����棫h��*>�9`v+�Mt�ļ�qH���q�(�(�|��1<�u�hs�3ZJ�J81�Q����X�7]�p��~9^$d����o<�Z��=���Д��Ţ��Z�ջ~A���������ꥹ��X4�&����'�)�[C�l��w�V�Y0�į�z�z�,$c�*y��B��L���@��1�=$�A,Qo^�D-�5$[t�05Xk1�Qх��5��ZĤ_�U����~&�ܴ��v��v��V���b)-�a�Y�?!�G�=�u�EK~��`|�@ˏ�����n����+��iE�_����|��!�r4�]Z�w��ț��߀z������<�(�aZ%`�Vj�3�U�8�N_y8`���̟?\1W'�����gJ��!B\��gZ��\����4�� ��E
���\?A\�<Q����]ǅ�+<Ʌ���fj*�	���6Ǽ�2.ܜ�Io�ul�\2�F�ǦD����V�t;��Z&6 �.3���S�G��#��fJ�����E����%��V���O
v��-^Ϟ�A�Z���XY�t�,���g�&ѻ@�'�,:OwC���E��Z�t���ޅDf����X|
�`J�{}���v;� C ���D)4�����������տ� w��L���zJ�.��C�vkɒ[Y�����d���^���^Ҹiѽ�kn��Q32Fu�<a�is5�	=vf=��@Q��m��kX[�	a`�.o��2.���WI��r���'�Qq����t����v0���&G�ڊ��aS���./s�-]���BY\B�W���<?�c�+�5�ԑro7�B]��~>�wlj�`�$�ɔ㶎�j`�EI�.��Y�ͺ�C'�� ��[�L��!��՚4%�y�"/]�Z̗\i�%a}i����\Y��<?���d�#��e���cґ�6ɧ񪃀�X;M�)����.f��L@��SO��,��5yl�-���ޱ�02��5{ƥt�x��,���̿E���E0�,	uh��_�l��=)�cAM���R�=Dd��L�����X��~�Sy�?�:R<K$1�Bu���9ܡ;���%�0��v�0b*MT3bP�o�A���M��HR��՛>k����`B�������J� KK]�[m�E;rD��c�F��{�s�=�]��ѽ��7�ռ�W�o��L�·w���kn�0�����D8��<�m�O�vv����b_�)�r�<�� ��cI6	1#�N^�=$Cj[8f�r�#�A d�����25٪Wѣ��>:����I�l����TG�B���e(�<�4��)���K�| �f���~�����ڑT�䫞D�3�z�6�,�0��7��0:@���[��.`m��>�{c�D=�K���ܗh^���V�WY�L3ɤ�έ�ON����w;�}v/���ݳ� ����#��*���¶��
��5��:A�7�B���˷x�*h&Sv+��T��O�zɳ�5��jϋ8�DG�HD�qxa<�E;C 88����N3�s��f���,����v`�(YQ]6��Soq��7��E%бh��>F�H�ʂ(;/�&b|�dy�YߦV�}
�h~;(Y��^㗪�B���m6�Q6U� � �A���zRS���1�5u�NC�sp&:��+�y���+=°���K��Ğ��hѯz�����6����a�o�[����f$�'���䩬�� ���^�x�;9{���F�m�@��1��&t�NJ!Y���)0���5�~�1݊�A�WC%�A%ԑ�-��:)p~ Z��@�����枏����D��'&����+�b�l�E|�G��K�؊tc�Z@�
e&|G:K�?�XE��){��)�sR�����Js�(�D�
����1�[�}5ڑ�=,<Ő����q�S���\�q��1C��K����O��z�z���Ox���R$=��;>)IA�q8��5��L��V,SO��f��ZB6�S�.��D��Aɏ����b%���펻%���o��(D��1�Es\����X胂�$MN��]5r��w�ե=������U$s��׳): ��Y`6HsY��m.���;�}�.����NKck�f��eQp��`4��[��
H������6���P��us�}��r3Q�Y���4�L��I���^�{m�j���[�#������\��e�g��`~U����:b�<ý��^6���R��k��Ӷ+9�>������N%��/�ψ��(���׶�k�����y�)Ȕ\[<YWq���jF��9���B�R�w��m���8C�}(v ?��HbJ��vp�ܦ:ԐY�������6Q�5���Z(ەn�:ݗ{4��A��?@:�W���ڡxҪ�^���B��6g�jr�jd��w��/k03��
��ṞwL��T@�h� �M��{��%V{�f,>=�J�p��0yR$�8�N��R邵�Q<�_p�P�Uؒ������X���<bHW4:��@�\o����zP��8<�B��f�ռ��>�/�����N��j��;⣵����Cz����H�o`%&����|}G��_!^'�`�!6Ւ����K(��Fg�|[!�J<~��D�"Rr�{ۋB|�W(�Pꓔ�R��]?{����WpՁ�
�9�+M���Q��3f���z��?��Ak:��2E�� �wC��&P[�"󲣞2葔�L���TF�u�@ِ �aC�g�t]�X�q��������.���c:�L�>b@�'�pK�9��S���%j�F`�1p��ZE�R^�p��l�o�P2�eg�"ʦa_r��b�cw���O����J�-x�I�=��.��y�52\�?�nYL��Dr�˧�
6>�5:zH�=��9�����S����W�/��S`�Kq|�*�tE�*ē�9�K�jn�iv���qڝ����h�u��/�痩�s��ޠ��⎪|AAg�;��Ħ�g�S哋<���x���xE��l̴��G��϶?�j�
#�����[�}m�c����G3,�A�n�78�' 0ە&����O�@�x�n��{��L��X�^��e�Q{�"�e{Ô]^����*93������u^�xB��m1��*�`����݁C7[g�!�gF�-���ë6C�a>�;7���1�/�o�ٽ�6���W�y�����(�Z.��>�U��6p��+Q��'�7��@$iT�>@o�2F
��U�moqc�Ԥ ���r�3Y7d��l����w������Q�ƙ:�l��NpY�3��5��.ư_wG Op#�:���0�dZ�x���F�D����rn׊�F�4J�vN��<mG�����/)a��훼{�w��v4�=6\Ч�h�jxss>�B�޹�T:+�k(��T��3��$x�����Ƈ&N���lx�0���:���D/k�4k&���]�d/�"�C�:L��s_�u�hr��ϭ��٫�z�R�#��t���f��#:�{p5.*�	J%1mx�����u_���6���4���o�g�?����D���Nŀ�i����P�(5<RR1V3M��0aD��Q���XR�

`��e.ּ6a�sy�4��ffY�WW���y�!�N̘y�fØ�;��d"�3�Q�+�OX��Ipj}��I��e�9���˹��~���`�+�2�i�\7�xͥ3���Y$?����K��UY�c�,�����f3�o5zN:��Z�X���wo�w�:r���/,��]mc���@��۳�ä�l5+�ʨ��\GZ��D�ecYD��/5k_V� |����-�k�}��1	� ��t��Q�N7��$YT��W ���6;��^i�:�`�B�����D̳�+�}���7����;ͬ�����JT�Q"�4lM~�~�fG��/p[#�Fj�-��ь#�$�o�%�?R�L�����T:�����7v��?�����<u�S���I���"�L�T�g���B��o{�"?�-�3+v�rs��<��Nߞ�&��y�M�z�D�K�l�/;Q���d-K�Z�4��Q�w�n��I�2mq��㝍����B�U*D/.0xY��v���9^���5W��Ţ���<����r>��7y\�|E7;�&�^x��:��& ����
>�F���2�(||+ab*1��"ꋃz}�T��)��p�׵����J�r"�f�cd�m�)��^����O�����5�Ҁ�>'}%��P�]��_�B�J��eci.VN� 2�mn��8�K������-�4�;+)�C�@��8�˚���QItjS	�s��z� O{�5:i�T�2:O�2"X�^�_�NR��-�QЩ2��AM=̶�����1+��7���q�1	��HuM#��X��B-�(e��G��|�����;nv�`9�Z������\�}P��c6�QMs�H��Z��u;T Dw��}N"x�A�7���Dd�!�2��[�C�[v���/�|5�9��3����Ug�y�< �~�:w�_���}��r�A���0>�`�\+���#��!RD�L�X&Ԭ�"~���R��"�h}-(j~�j�j2���:�DA+W��ί�'��N�M�
]mh�P$�@q	Nu��#ĕ�����]�{�����r'�w�\�!4��Y{A,�6$��:��ar\��xIp���5�6`E��ݩ9���t븖I9����r�	E|�j�,�jl��.���fߌ��u�}.�]`�u���x��YYㄶ�w1 z.5)�b��Y�t��:��hUJ�C�a��ݑoGZY=�Ι����h��噜�
����(�閏y(
��*q��_ħ�gË�2��h�=n�|7u�u�p���N�Y��tJ� i�v/��s��(C�7��ȾfI�(����V��rM�!������5�TH��f6�ҏ@a���fR9���K�^�e);ǁM��B�ڻ�1x�eك$�9�)&r��	U�$XXP F�w�5�O�T��VX �Y�t�]|���'���VR��y�¸�*�`7QP�@�#\�&a���M��n�� �G��bؽ#��/UU�h�
��Ey�Q�]�q���튾k�9�qX}���#�A4�V'���Hi� ��S�����V)?	�e�X��	��KVJ'��ȿ8�l�1(�,�.�ًM'k@���N !n�^1Ѣ�%�_(i���\d��H7|/A7����]�\�hЧ���9QqZ-�7#���q��S�?���"?�9?�&V����xy, ��LW3�r<B�,�Q(�Kk4���� ݑS�E�o��D�0�O0�J�� �f���uŉ����,� Hڱ>�t/
�ʥ�Mg<�2=����� 9,UK��cB	�$`��EYkFiH�
�
�P����??]�Z��-�
���I#�hZo�>@��`�����t^E�3�	!*ɷ3�p�(<"G�ځ��R�"K�7_1�#��}p��^z݆� �"�_����&}��ݞQ|`d�E �ݞ	��ߘ�s��z���=�5��s����nr�	=���$�)���?�/�P�5r�m�ax�H҇�g�;�]x1T�+&��'���MR�(R�c`g*����59�7b�E��?�#Pe�Po�%�:�| �D��F�t�e��?)�kC����m��O���^:Z���Q��?��'�t_�O#��I'h+p��u!Y���4N��#���wũ���i"0��R�#R��t����*'��h���S�h��"�����{��K�:D����|v1�thI�;�1NȀ�-p��s���W�����U�4W�<$��h�k�="��>�� �Lv?ĴX���8}G�aė5�� K�b�"�ό�:Bk(� ��w�0����>����º�J�ƪ���<尀:j �!�/(+�7���+��9��IP��Ơ6�G�d�/�&��S�ׇ:YtAE8dU2nBp��_���I�o�G��0Y>���]ߣ#����K����h�-�<e,pG`��cM�ՙ��k��S4۝ޞ�Y$������O�J͟f����Fd'�Yjg��'�(�b���5 O�(0y�O�9,��:�9ڹ�J�w���ț���x��O��H�-F}����
T��=�)t~V��0�R�qĢ��5�Ыn$�&f���>��uԩ�F �з��+"��T�ܟ=�����yD=�S~	�&6u�&l�4I���5���_���ǫ�2s��F��Kק������j�!B�������?�9]��D�JJ`?���G<�V�I?���({�χ:+W,︪'�l	�Y�5M�ϵ�mX�.0I�m-'�x��&>�tg�3b?{������>5���|�J�U~F�Jҟ��| �m)�2�YZ%|�3��5��Ks�V���a
�a�Z��v�@��?i���GWC�yS�/`�Z�K��ad��8�W�";ߟ��
��� �+�C�cgFkD,�&��ߏ�p�{�T���_J� ��5�{�Ym�@ު�Q��oN�{y��c%gblQ���H���ݎ� �فQ@��R�y'ps���X��$�Q�Z����ֿ�i�R�O�kޗ�=h�°��/3�Z���x��8�,�N������Q���ߔK٢�(��]�Qs���5Ǵڶ�+���S[���N�3��U���=��n�qp������-���P���Cu%<z6�l8|��c���1O÷��@b��ma��X�L�e������Qy�01�T�����3T�	V�rQ�m)���4~�B|�n��a,�Ќ8\�D���8�B�XM��l����*��s_�sm����3m^^��C�V��w�����b`JQ�0��ɢ�}� � 7�l��<EW5����3���Y'��R�\&Լ(u>/����jB�lÕf�G��G�3+ܠ��t1Ҩ	��r���$���z��1�g��vz�H��r���<��*�\��i��ӑA �Nb�Yz��G|�Ss�܇ڶC��F`g��oy�ԣ�^�g'�	K�uא�cy^XM���be��c�Q���Wo
��D"������d�j>3'�kC[ç�9Blu����� ����+70��~���f�ܤ��:�-|Nw�7�X�4�P�8:����㪠u9gn����;��������!�x#t��OM=�����K�}��@'G~>��	 �u��j����g-�A`����=�oE�m~���&����,F��\ݽ\��zQpg�b����}Ḝ?H�^�_����oC�l�Gz�G�v�[�3��PF�V=RD+�+�/_�Hh:d�&����G_C�*v]v�o�Fbݱ�<Jk"��A�P�N�|��u!a�:\Tqe#��S�}E��S�Y�qO�Fs�?/�����Հ3�U�>_Yt����D(U�G�_/�D0pP���;oJ������{�g5��`Y�]t����om��g��Ɔb�C;��X�N�"M��2m�m̙��cu�aA���@��������"�"x��c�o��p�޲kn��UL�B揤J7��S�Z��*�,�kط�Yr�wK2!²��� �	��%��d�Z�]��o}���2Y�c�d��8uɸ֮X�sN��]S�V�ld~c�x�m� ��N�yS�ib�e��h��0Z�	=|���*�����.�`�L���Y�X����6���y��P�	P<�}|
�#c�+��Y;u
b��B���*H�)�s�I�1�?q2r���W5q�`�� ���Cr/	���#ۋ$@���D���1+a�ۚU�~U(#B��ع�j�H�q$���u�G����/_���Ԗ���K5�GFMR�z����o�l�M��A�!R'���/�`��Zc����	l65��������"E;�B;Gq9<R�2�G;�T杻�W=a����?F�����g�@16���K�J-AW ��B���S�b��S�����_ی9���W�C65#�!��3��b`ެS�$�T����묊�Z��F-�P�!VLQ�^�0`C��ѵ�E���z�+�G���`�K� M���:�g���iP�b6�c�'�d��3��y?��i����
|����Oau��϶T�j��C��X٫�r��d�L�'0�k�����<�YI7�I���ܒBZ۔�S�f���
X�+���j�lضDK&����ɕɆ��?��oi;5�����m�o�-����qZ4C�Jt���=�!j3�4�W���s)�W��׶���@��"�pŨ63e�h'hTi#ҎQ���;鑻��f8���=�f��ot|3D����C��[<�à���
�[`�����~Հ*�?��u>��Mjs�����Y�wx�R6� �t�п��-4��v���W�[�����eg������ۋWb��N�(7��"�U��+�����w�����͹n��Z�v���$����ޘ�{��rN�|(�vc,���)+�EVoJ�F���]TB$ъ��� e�I��^�/ұ�
,X�꒖�6�����%	pb�ȶ
}S�	[��.�gl�B��P� ��P/��a��w��8�0O�_�<�A�C4��a	Mܜ��qc��.؞�s-�k��D'KE��pAh�{^=QA��T�}ȆN}�,}O�m|������#���ek2�o�y�+3F�E	��L�Ѩ�<��A"?z/��lE��/���tN�u���
�]+��>�&^QF���춣��};" ��ܤ��萓�]��b^ Դ:�c�zU:g�����wo��k�o��_3�Q#2
�W^����}B^Sg.O�����t2���Dd��.B��_�'�ޝK����G�2��޹>j>�m�FR��H�sL�����ݯW_�`��a�e��	GN����1�c��>(��o�'u���k��}�d7[���_F��KaN�����J�r-�U��\\��9��nѦf���g"��0D��Z���c,�i�e�UO�j��n��h\��&y���G���P���=�Sċ���J����l�Vf����6�=�7��Dt���sC
��!�N*���h��:; "��/<�2�/o��U\�17�#�F�#��`s-�`�Gg��q/ç��#Qp���#��L��;9q����"_ͭ�J���L�
xa��$�b�!{Ҥ���rys�_,��%<O�Cm[b�iFuK��@���0u��^4�m�����:&��al�<ȾjsѿHI`�^=em�u�th������uN������U`��X���e��ޟ�ʸ<��pP��Wc�tK�,n�Woi�,�����Q�}�����W��\j���;]M@�e�N�~g+<�k4%����G���y�X��]W�v	 �z�Z�w3jK����g�-L;��G���#�s�e��#K��d�A[���+`�*�Qo��W�}?ZG�BJ=2��V��u�3M''Z�k���-ߧ�א}�����	��Q�:tQkk�8�A�9�q�P���!�٫��r�L�����z�qfɮ;�󰸭H4?F����g�� �L�>?�'/�������{�ΐ�z��Y�,�ጰ���L.z�|��I拇�\���ćE�4�w�=�a���A�^Q��X�j��.��{7�Nqӥ���;װZf����.��&�rR�'�������AƐNc�J�͔O!\I�7��s�B#N)JA������֭��أ4���p�-F�c��$i���xRZf�"e��5t*\�T5e��I�Կk}c8�d`{4`3�-�q9���vMy��{��4}���U\N�����D��yt����j);�$�\-�684[�>���3���+���<�KY�#�d' ���܋+n�}�~�Y��-�f��(�\ՠcݬ��Df(�� F�"�d�0,٘��Sm���
���k<�;�pCjN�.���9:�=�Ar�6eqK���qt*�{2��|8e򬵵&3��cdn-Y����Ƥ���Jv�z'��Qy~��ebI�;<P9�����ⶼ�,|P���n~�7+��}�Β�a�4�zPd¸g��/Ɔ@�OI�|a���E3��8�p7%�f��c�!�"8����AR�����05Қ�����{�]lG���j�i7��p.�[x��!�F�eN[�s.�a�v+8OP�����,�:�
S	��#��z���DϘ�ȂN��-$Y����OJ�T4���v=lAo��WH�%x�^yd8����q;*ݫ�,"\�����N�����D�z��EL�E��o�
��P�=�u�1��Z�y<�I)��9��N/'}R��@�Y�Xr.^�9|�#�[m��|�}�u2(�떸Xb,���T{�᫦8	��i��ź�P�y�%�/�A�pv�̲�d�_��T�p���S�BjlVllǷ�D�^����� �\7,{� �믰��Ӫi	3�
��y-�N7��%�z=B̝��6��2
N����Uh�:����ᯖ�M�J{��nBT��|�D�K3�b�P"�#O���7�zV宖�M��k%v��A,Tح�u�F�Y^9�h>�7R+�6>��YR�~cN"ġ8��.A&i�\G+JV0��'�1�I�ᕜ�����pX�bp����� �$�1�j����p�$��S+�������,F��T�^�N�g�l�Ј��,H<6�p����9i�$�N��;��%���^&M���j����4#����'�.h����U)w�#�f�%�e�Hk���sB����d���.�C�U�?������{)Ab΅��D�������/xx���\s��ڹi.�B�: ���U���1X�V�fS�u��\�
�lds1'+,��=c�m�Y���k/qN�fB��	�6Y�h�'���l}�{�n�#�5GB�j�~����pC����u��'%4��fk'>�W�{���_�cfUI�Yv�d�]��rw�
�RW��_�܈�r�����w�{��J�{hN�nv�O��6b�ڄɒm��ѓ�p��J7ʦ;�'p�n�b:t���$������a9��~{��w6jo��<(_�R�sȐg>m�h��#���m���A�bl�z��)�磦&�8����K��=�����2<�-`R�%Bf�ٛG����}������\�m�f1�L�x��t��G�y�C9�qSl���KZ3,�I�	E{�i�`��u�=��`A_�mGG}�{&c��_rCgv^��6��f�P�!�Vʊ5L��n�/�~Ͼ�=j�z���ɻ��\yvR�Zf#���z��:�Q7,��j��њ��8|xI	L�}G�n�u�7�e�H�x�sq�"�/�^ėoU�RG�;)�F利B�Kq��o��?lʲ���ڢ����WLxDVNu3��>��g[��I���
��9L'��-�[>Af��u@ZS�����W��*��w*0��������)oYY���iX֭zl%�"J�u��Ts��~�a.�����k�AوpZ���΋Ǡ����hc�Q��H��MY�ĵ�ױH�����_qD�p(h.a�嘡�v�_�S�����YA9�s}���J!cG�!�b'^� ��>��������MMϦ��!�Pw�����o�{�W�:�\!��'�(�j��6��8���\q����A�P��K?��9���Ə������f�B48���������&��M?��13���W�Ӿ�ut�2�Ў΀J�W��Wҷ�xF��І3�!m�V��J�I��f�M	�Џf�W6�oj�1�gں�cn�\�4�栾��.����G��0b%~�? +8배U()	���6��jP�<�K�������fsp�vz�^��ς���͗�>�߆��./{8~������C�)�Ad2�ٗ���Y(〈��v��T��-�G�"��g�5��b&1C���cm��3i���5s�؁B��	AB����@!�1�yJko�v(�����I٠Sr�E����^�3>��U��} �=��U�E�͌�&W<�rKL��w�tSI>5(�VĬ5T4	}c��"r�z�}������Pg�YLf�X̘Sr���_p�ɴ	�q���N���p��;S�^2EƬ��)9�M����ܱ�13X�P�zߢ�+����E�]I���8��5^��Q�69�z�
*���/1�)a�}�Vd��w������lt��e�E�iw	����6c���B=�V�$���:�Gv��ǈMΨD��:��j�p�є���k����>���F��R��h�n��V�OÑ�vk�Ay�8Y��ͣ�r���L�b5#]���.������>7�������sM:79>UiAlN����-���8Ư�e�+���2��Q�$��R�U���?����.����5�m8�9LWF��T1�[�ʎy�, �� ����Zٱ���꺔��"s��g��Tu�xw-] ���f���75������|���GLl�# �<��9v-W��Xg�H;�׋�Nl�S�F!e}����XN8wle<˖j��xt ��+�����=pZ��i�?�3�x���2��~�>G�q<��0)}�'��@9�VW#��P#C��,�d��)���מ��ѬP�����ݛ�փeT�����Q��5�Sm���|�7Ψ� lуC��lQ'u�\�:._�+��NA6�5����Z��I��wy�٣������5ɋm�ۂ��k���{V�?^����h�e=�P��E4/i�-C!��f�t=L�+԰c��>U��4[ǂ��EC	�)�|2%�NK*'Z$^w�4t%�V�mʣ,έ|�x&>Ǔ�r-�7&cz���jjF-X����f�3��"w�`a��@ �N>`�e�i��ώ̖6z֓�O�i	㗚�>Ry
'R��]��n�U���_�9�:,n	s&F��Y9c 1��7#�Eds؁-���T�o�Щ\���f��p �������i�>NL���*�5]������v�ݒ�������X��Ӷ���
�����_ݨK�N��R�տ�V�*�f�[t.+]iJMii�� 5�W?�wh�}u(#O�O�}m蘙8g;;Nen��R���z>tW�����I˯��#��[B_�������g�7PR�񐁫C�
�覟߄�p�$V���YπI�cN�l�Dk�m�Dɼh��;	d?�1Zp�Y �y:23�V��w��8#��O����`^x	��g��/8��ܑ���J�c�*#m�]kV+-}'k����q@p춁h8�p�v�.4(Q�ۼ��6ۍ��`��(��&J1�_�G �7lr��͛m�)H�M�G��V��E�!e]���~�W�)Γ�v��4'P��P�+2>	F�w��=����A�`NL�$4��y�I�<�4!��^���ܗ[Ss�G �m������������uQ���>���_�k��ǖ|���Ό�����DdI�mߛ���Ř4~/�s3ҡ��D�Uu��ġ������-�̸��web
~����&<%:��;�;���3�it*���?q��;f$�J��}}���x��������O�֤¼s,"9�����ȗC�lpڲ�7T�Õ��YsȬ]>�Nfoxm����¬�G��}1�ۊI��_Z�H�	63
���9N��yY����G�~:��y@ݗ:e�eՎ�����%�=+���'ԈHw[�f��P�J(�jl��@+�_0R@����T�!:o���p��H�����ǺM�)ߥKW+��(�R�,BY:�>2���p�J׉N�`A�Jf�� `i-m�Z&'k-���|����l>ӝ9iQ-�Ժ��h�	�g,�	\����:WI�߯�s�|\�����\��5h�vurw"`�Z�ʌg�y��e@����`�-�@0��������(t0uHt�,#u�F�-��/n�ڜ$�ˌLO�������k�^����x����k"�&�.�a%/Q�1� $��c�l����5=2c����ed���2�#.J�I�c19#�S�݁��8�(�8��c�dN�m�Q�WyΈ��Ú��0�Λ�{�j2EK�a�T,P�KH��u*{L�L��S��q���t�2���D� ���R���C�Y�+b�+U@�`U����b�+kO���D�X~�!D$��x�Cy��ᬷ܀�[�W�S���� &4Kvz�L-�q����[�A_�M���{]B0z���, -�X�f�����������7U�9d5��F
G��R�D�����E���gk�9��!2s	��?�Z]�gȨ���D'���v"n��pm��S���,Fo�P�ix�� ��+/�șu�/�tL�r��İh-F��w>���%����� �"���?�?x-�hF[�|q~s.G�V����բ�!�\W,�S�V�Z1ܑk>�{��v����P!2|�	~��̊1��n�f(l�*"Ӷ`�[��[=>H����A����׊=�����'w)�?\�+�}6;�_����y�	u[�z�u����fư����C���c�� $�B��lxg���{�ow����S����(v�ȉ0&�ΝX�J�ލ[�8A�R�ü��ͷP/� ���2j++=`��������I�����wl±�U��p�Z�*��芏��J�����Y������)0١ϩ��b@�Z��M��a:�ޠ�YRw�r1��)��0�#����:=ˑ=���~�!p�*[��|o�:7󾗞j3�(Jm�~��с���'���Jǵ���ND�c
M2+���F�Lh�`���&���,�����S��<���~��^�%�q�l���*l��!Jf�D���(dI֌^J���OdeE�W��lD���"��˺wsc�vf����g�t����!Fg�B �7�:ϋ��U�W�if���
����؋�u�G<癅��RC`�&"��
��[��+���k]>||�F,4�nS�� �K} ��{!$������!����AA&YTWV��M��J#�]�x�D�b<m�%ۭ�%A�ĕͬ��ß/8#JQC��u"�/<��?]����KF6�a��)Y�N_*䍶��������2$�#7r�q��vc�7z�V���=sG��6��aI�<14�~6�����#1�ס���	�B���UM�BT����T�+g��J�!y%/�\�8.���Lv�"/��2`��|�9~XQ �4�b��ݟf�]/�c̙�O�t�h�G3Kz9�2m:)�}>�s�?���T� ���=T,��|�	�^J�A�'ˊB<0M��\{����"�Tb�g�=A-��y�Ya�;Oi��@F��ᙌq���F�YQz<���<���7{�j��KW�x���O&�Nq�Փ���M�y�\ ��J��ل�Aw͐���ڵ��0�O�*_��6lg=/r9� u�S�/Q�-<[��dsz' 4�W�')G�ɣB091�B`v`����'VP6��$��|ՠ5$������(�Y�F�������L��\�f7��=�^��48ȕ���o ���,&���Ŝt��I�6��=�L�;I�R�DB� � ŷ�L���9w���E��s�q�a���=����Ӕ"F���iW���s4>?��9̬H�4������_>���e]s9=��q�)��rJ�f?cX�)GBcOJ�<�����տ�:����
����9ӏV�ۤTIiYM���{QV�;��L,�Ue�* ��t��4%�)��O����5A��RV̼�%zZI�K<S?��̓Hd�MB�HcV�?p��9���M��Յ��'�8��!�c�.������=�y
qTև/�]��&������8#b�͞�n=��bS��t��R���V�iۢ��d�� ��dF8�(�D�>?�x��+�����k����,�}�9zB�X�c�72m�zSN�s��|��.k�-B�"��(�[v�$a�����X޴��҄������3�d˧��	H*���me+�"y��U'ħNtZ�9-���W;��겖�qL/���D�Y=vӽ�㼬�EE��6����1�d�B���Gz��F{��L�e�"w�L҇tj� &���L9 �h��聡�'-�7�c�6�-�)�- CY9����so�$�5E{&˞g��w��X`�b�M$��ߤ���,�x�x!Bh����_17�3*_C��\ ���DF�Ŷ�o���:�v� �d�S֩�m/NU��2ء#�y̺|s�+~��� �UO����[wԾ���ɡ���Ω8���~S@Oi~B���ެS�NqFي��|?.��_�7��F�(��Ǥ�hD�% �c0{a�݃�� ��n�]�e\pϾ���&�|��	�]/�� >�_�5hH�E�*��F㪊���f��~���U��'JҵM0�#���lp.��w�%�
�
+�K�d s�g�7��8�oVn���b��_��t�~��:�(q>�x�����}@���SME]��M]��������� Eц�ݮ�o{"�����~�5����r�e��s��R�5��쇬�ַ0�F�{e��?@4�O"􇵗L��c�E!��
&��;�/���諧������,�_�y��?�}�s�u�4���yOi��f��f�܌hq�~�=��S���K�N�dPI�K�A���'� ^��L���+��a���e�kƞ��ؙ�r/I3B6�����t- +��:��5&�s�ŞA��ܓ(�;ez�A���"e2����l�H�^�!7z1g�ҕ��fϺMʵH�XjD��\�f{�z`�C�2��
�3�Scf�7�8�lI�Z�ur�"稶�ǜ��v�{ԟQ��b�
(@�NE��{0`7��IJr�ӡTIz]ʘv՟y���=J�U&��� i�����Z��>NC�[���kJ����ر]��HyZ�UĠ	h��9����0��4�*��q�@�8�PW�ܩ�J�����؁����+Ao��w�!�0��:�tK��`������ڳ�;u�)�p¨���,�[���	�]ELZek~�6�_���q�}�G�z&�h�"�Ř����j)��a�v�;���4�[�-�е7[kzGbB��%��j
��X&��^a2흘,��dv?�?@�Wiy�r�i��G��"�s��n�=�F�}ZEP�,�M�6q���[ގusIv�+���L�j��a����<�R#9��i�n��K]��Ù�3�"xLT�ȍ���>���-ܽs�/�2���@����P�Nޤ�Ѿ��%�L<�dʘo�.���$������G�μ�!�����T�Jx0����s��4�L�S}�w˶��X/ojӽ� 0�k�4p S�r����ֵ�!7��U�E_�u��>�+qef�{FN�0���s��w�]($<���D�ۓ��/���W��G��'1*�e~T�|vO��+��j>ԯT#H�^���G����DJ���4Q�l��6�~�V�%������ ��Q!�]A?�zx��Ko*�H~��*���4�{��V�M�G�ù[��^3��K�;�Y[�(�l�%�L���^ʣl�"��d�i�������@#<D]xc��Ѣ�.w�L�E1=ۗ�}�XMU��&�mVt+�BZv�X)�����ֽ>alǾ���t矔�I����З ��µ�������.��5(�&&��z�1Zwq�U���.��xi�IVnO2��'l!r���M�[�G4����D	3
�OFG�,��Mhp/<�]�>JM��K�Oп��E�C���I[<�@ު��jël+�{�Jw�b��^�t�f���7�G��	�*��o�GO	�����m�Ȃ����E�P��#k�c����K7�����XB���|'�~�h��j���B*�]����%t��x�p����F(Tv�B��/n�o�1�˗����7u�ȫ=�1��sf�É�����ˢʅ�ߍɿ,���Ǘ�T)�����4���#��L����F�����#+�#0Y�/κEAi��A�5ϔ_>|��|Q� �J��ca�������T!6Oc�*�<�2����Y��b�1( �RZS���I�Ӎ�Jڼ�f�K��v��]ŏ�^pu�Á���ӛ�S*1yC�,@w����
��[��� 1�9\j���ܪ��V�Ӈ̷a�UEB2{u�v?4p�.oq���38�>/UI\E<�'
唙�K� �ݳ��Qa"�F��@�WLa9�t�߉�H��J�h��zM��ozʑY��m�bH��w����M�����8�y�%��QM��ǈ�9�`�I�Ǩ)�Mݩ ů���H�	,	)x�z���od�б��/	�Eހ��/���~�L���
��/���>��Ӓ�M���M�Fv�%��nWp���8-�HC��;�C盗92��'�)�G�Vy�������CQN@�� ���YV��aQ*.`ʀ�~P� �,4�A��aNu�#	,\����N��	
�����W!{ �<�Uz"\��N�(�K{�cyl��β��z�y8��U��\�ҩ��b�4� ���u�JS���p�H(	N��T::�k��r��s;kt[�ui� JӜ�XӸ��M�ɫ�E�[��4�4X{�]�`��{�#�貳����h����Hڋ2��8(L���!��*#��m�Ո���'��2�2 ��<���i�S�s�:�Z^�d����5za�G@�_�x���ܸ�~�hP����߲�������C�>��Յ����s�fro�>�
����:�+���i�A\����n�Y�%,��mk�&J�Y�sx���(�������Z��[=���loLI>��ˉ$=�	�<`&�0Je}|r8���Y�	�Hs���o�tSb*;'�$8V�7l
�g�-j��5��_&8P����0����Xz=ǌ�]�H�5������agz_R�u=n�@A禙?;��ֿ��eQ..��MN:Jy�!��6rtV�=�x�@�nA�#p|5����2�`@<��������٬psm�M��M�ޙ�J�%����4����N��d���]�iUI�
+�h���ڧz���-�^��y�ʣ��Z���e��jʍhF�{x���2���F �]���G�n���V]�LL�BQ�3��RC	%��%��_�����*��c'�o�Y���)�07���H�s0������_ ��	����}�Y-���\�#��탹��B�ck�����,j�ɘ��4�`n�-���}��Y U�b���X����fa��`q���T&��7ᆜ���~fe>�]���):.}!0@x�JC|h]�ҪO���(�#5��Ew �.��þ՞:(!��a���g�N��4C��]��D�c=����RO�=�A�ʇ����H2x2���O�˴|)����qKc~R�1�5��^5�2n�űHk���s"�00�)��'�ރmx�������d� z�pV�XB�V"]�6��-�HX��J_�,���uܤ�zW��m�ܣ%��R�'�L�h��(6���k8�����Uh�CK٨;2HY��}qA����ę�ב/�Ş��LHOX�c�z�N���ަ��9	aA֫��m2����q�d����Y�s ��`)��HuyD c�J��!w��	���xI>���J!E�Z`=�*b�C���x*�d��ʳQ>��H����9��ٸ6�8}�!p��������<�	IZ@g��ƾ�}֏���J
2�a�n Y�+�8-�E�.�΢��2 ��\����t��s�D@��� ?S�#��lt$���M��P=Z��o�ȱ�i��=#̕�.%")Q dD'�an���_z�$m���w��N�J�pW�@�8,�0i��k��Hгf��_��ol�!M�9)3�:��H �n?�4���q
0`NY�s`)�M�g6� ���ٖu�o��n>q���J��	� .���� h1E�傤}4���"��a��qM�n �̠�� �s�"��vC3���rpl��r�[@�0F`���:�y����x2[*A�u!Q9��n�J����;�J��dno.vD1�wS���7^=8���#biT��л�Ikx�p&�FL�Ǩ�{v�=[�sS��U�*Ӂ2��(�u�o��E�H\^�Ė�U�a�E�&�8ӑg��F�5'��q�R���K����l�/C�pGV��G��󗸬���Q	�=ϗ#�tOenIi����ܿ]�f��K�/X� 
/�����5yU��yH����p���y�B5�U�v�zq4X�?sH���V.�:�M��6�q�,;�!E����? ��8�	�;xo;s�lZ�7�{u�
~�뷅G�&ܮ���2a�zQD7Q9��/�O���&��^!�@�(avA���u,��/ؑ�}q�
V������Uɞ��QK�v3��z��|��h���x�~\�22��k�q�-�I��f�#����8x0�՞^Ɛ��
˛Pv��SyB�H;��߳�\p�x57�#�S�5�Fz��w��R�����<	{D����K����m�����=���`�C�	�Lr��U3���W�c��0&7�:;�$jf�\�G`[���}��|���On�����l��[xr!��n��ε�2�^���z秝���]��K��TR��AD�d�3%=�iV}��n�^�Q���I����0�<᝜L��$꧜���:6�2�(e�֖C�k����*u>�u��؈�Յx�-\�����w ��o$.�q�~�Y�sO�&�1��,�s��&ք˲}] FELc�����H�({Lh�)3��D�C;&A�g���j�S�9=�?�����f�J�N�E ��/]��$^A��5e�����e��d@Z���z ���+��Qy�g�����{��Yr��s��e�=߿R���M݄O�wgaLCn��v�ᡱ^�X��3�����
;D2�Nt�^Ot��=�2u�&�9e"J �#wuV���-)�TJ��i��ܮ����`��ʇRWaG�t|�0��N�|ǌ�t��<!��4��Β"��иh�ҹ��,�#v�T蹵��{�0Z�H�b���[�ɯe���ɫ��{�S�t\f��̬��Tuk�O�t��{�T �6�k=ޚ�S�����d�H���KQ����;�*�V(�츥D��}Q��v ߨ@�LF�����`��nL#$Wu����j�}���q�K��y�3����3�l�{[�M&e���&|/$�j��m��|���v{�d>g'p.��M�IX�ڦ�$d��:�if�b.�fz��wK'�,����;[)�v��Sj�&ͫgyĝF�<D%�5^��:��*���q�w{'Ѻ@�͙��@	K�0�[^ꠌ����2xkp�%ұ�ߺ@dS5�^�@�/�v�t#z�/5�R�hǡ6�KJ��vy<��g���N}�S�M��/N�G3T���B�����՞���E����� A�5���LF�O��}g`/Bt�s��^���Q�1}c�82ڮ���� �|�c�R+��1��t�N�]����V�`��^�t����L�U���w�cLNd_o�IDm&������0n�y�:���kbRu��:��E�;R�8���_�0��Ĕ�(Kw�C_�]�>O�y�S�j⭖V��$�w��oR��W;b�s��Up���w�%6%9Hu�k������	Q+j�c��p��S�u*��9߮2�H�a�<}q*��Qh&�a��Z��w�s"���"ҫT�:�v�,M`f�$. ����P1k�P�꣏�&�>
�j��H|-��@�!#Cg�~Fsl/��@^?[���k֒��3��&�?�m�~�Po	��"�)��2������l��~���i�b-������OJ"������Y+l�NO�A�Ď^n4W=�EׁS���R�1��p�[���1$���7�����aB;���t�e2��4!��m ��N�H0�Pw��֢b#�_�N*�M���L$��&u��s	��.�/-��g�Z�A�|�;��Y����|*��`���nu���WGp	�/x�ƒ��G�#2^�Q��, 5���K����M�`�p֪>(L&R�>���^��>@C��`P�(�!�:O5�秙�zֻ�b������U@�����{.��iX��HG�כ	��_&�3�AiU(��tt����_���4"�^��e8jA�t>	�J[���by���mˀ ��͙%Ź�Q�4�A}��7Ѥ�p�z���Hę�_PA����y�fw�>r;�����J�^an�CБmb J�
��aL�]0�ZQz��4����B�+.��P���Ò�o쌅,��`ZF�<��u�>�������f�3����G���<�Zd����y`���J-&�\��h�|]��l(�m��[�5ҋ�%��F������J�q
�
ɥ���+��hL�ڂ,��]*��Vh37�On���+Q�0�P�i�СRinȧ�����=Z1�`�^-e�6�=<"�����h���5�w� ��_c�o�����F1xQc�'y�(\p�v��(�R�.j����-IxcW��jo���^&d�5��t���#���CU�e2�DY%�͝`*'�~a`ܱ�k��y5Q���`�-�PI���
������^z�G2���<o��H`����{�])�'PEf�Yl~l>��ꉤ+��D�f2.�tB�'��ʭ�#������_�lu���8v�C�|�1���-�����Luu��P���OJ�W6Ǟpdl2Ү�N'<�O~��=Z��.�45Wl�/]�8�|����ć��Q܍�
��)������)�03�i]$mr�;8��ꖸY��[�i I�M����QF}&��������4����Tu��vc�b�Ux_:�hZe�5�༼�T�=��f,����z&'SM�(ՅI����!��|�L^��ϒ�ݴQK�����)�j! k�츅`�94~l��̘��@F��pQW����Wɶr��'� � ��%��fM#w�!A��Qe"��m�.�)�y�#Y��, ���ē�qF�̍#=&tvY�d�}�O��}�Uoil��~�N��#�K����9D��JY�qÕ@�l���f�I)U��`jؘ���'��Ʈ� Z����}ݗ<�!$S�VrҪ�Wؕc�:20b�%�[�0�*�({d�}�b���SF��y8��~2+@-+D/��t%�)���Nj����f��C-��J�]s̓q7��:�;����$E�g�����R�g��b����=@�Һ�шTR~�+���)�^�Ϭ��h�R����Dd:`�/�[��{�4����i�My�b��Q��[���u>�J��XH=W!V�Ѣ����¸;-^ֈ�֧K�XN�����w��*��S�>��6M�C@�iF}0�t�e���_Z�څx2S�6�OэH'�z
���W0���_�`��*m=Y��%?�#æ�l�8k�����a}�g0v�^����ԕ3��f=�j�QH[�~r�a3��yp����%�IR��3mrP�e�S�����!�(lą@�8�?㎈��0s+�� ����{��b���<ᦻ��%���[���	�ϙ�:D��%��{b;H��;��En�+�����"y�C=��.�B �����p�Z,���';+�eMq�:��V�.uk3�^�b�L�E�*��'����]?�q�&
�`O���ڠ����f�-�_9�~]�D�'�x�n4LH�y%E5�8Ү���?Iھ@�{�lQ
ʡ ���+��~�l^=�k�-���1_BW�@v�X�{2ae"ƽ�j��q2UϚ�ЧU��z۱@�ңk�s��\B���r�q^H�,�
n����cr���q�`g�]��]I���o��v#K���|Y����<ֹpE޸�~l|,�yʺ��{0!�ʐ���2�����q�].���6�{Ѱ�MW��E��7B�t�A�GF��p�$ä@qa�k�&���6��N}�`¬�^$�$z�����\9"+Wn﨓��>!��!�?8%p�ȿl��k�s|j�r�
X��JP8�E=�K����lV���lm m4j������(c����ib�13��k�#9,��-z�}��A����&�=mbҺ���%������eD�S�nÂ�Z�E"b���
+��ɸ饍�c��j�;hO(�xd-��	�$�)�4V|��7�ov�I�R���V����Iv��J���>Kh�Qp�ñ��Z��jW9���� Q�@ǘ��TR�{q���k��yL� �i��ƲI�	��2x��E�ʶ��H�����������?�����at�%��=	��7}U�a�)Ų���Z�2�9�@1�������u�S�n`���W=V�d�a�/��O�%2O��B֬9�R�.^W[<��v�{�ة��$]�]��VM'��8�g+�ߊ�`U��s#i���P�Y̌q�b���=���)��Vy3���Ud�_�q���6̊n�r2jV�U.i�yN�&Ԟ]3.�0���� ��$�~lI=6���pl{5͟��i%iK�-J�T���z�T2r�W�fQ��<�Q�Bai);�b3�-�4�o�ض���� .א�,'B�H���J @�^�Ś��<2@���O=q���K�?�]L <��Լ `�jx~�tv�� k���_����s���x��k�+���[�c~ ��SLw8� �D�PJ.�G�@&��sV� Z�FU�&{oij���喾�>U���0�Q�o6�����<Sv$��h���k\Y���`������d�����9������t�N���M�B���oْ7>lb���PJ����w�m�i��Bj5k�I����N>8�����41K}�;Hj���Z�����U�I=���7�v�V�0�@� ��kAvو���K��b�-],0l�ɖ���8���k���z�s�Y2�n���3Y�9�\]�i��خ��B���s>�/`��*�ۉhX}��Zri751<�nk�ih���̵
3�V�a�w5
���7���݌5�jS9�$���{�7�Z���
�b�*ɖ �ѠB��^T�b�I`f�Q��(m�9��8���f:���1�����	��a����s��a���F2J?>s�:�*�ql�К�r�`���=���Y�Nf�%n��N
׊�Ĕ�|�e��wWM��zg��`<zpI�&`oO��U�<eu�vb���p�GA1-�$�Ic���P2xH����n�]�U�sk����X����螀�L�KZy0b���YZFs��ٳ����.B�<2g��x\��M�ө# 8p<v����*x1����'�1��zs���>뎛q⾿��`�׭"z��!ٛ~iJ�����
�(@�1󼆃�u������i�gL)���iٍ���HF�4�����s�s�KQ\����0�A:�<�z�U���BL�K�)�߰�[�M�O�WͩZ�p��h}U7?�
3�@�[c��l~9)V&�)3'=�Ou���ѯ^b(o`�i��W
kᴗ@��g��.H�|�xLj�B"3��8�Js�ZԤ��COݺ(�N1�ӆP=@i�C�Y��2U�JZJp��z�p�a�mєd�}��;��m����b*;�������тKi�k����0/J�V��Z�tu���~7rB@�Zv�i��a�c?�m۟\t�' 3[�$R�[!Rc���}�dⲝy���nC��Ү�,C��TM|�ǹm����W�W`�8k������졲H)�w�O��{�h7`vef��A޵{V�x�O�]�]��
)`W�k'�f�e�T���Ҏ��sׄ���)��D�IG��
)�
	���^M���*}Ƨ�`C�=����V�a�T�l�զ��Px��$G}�R� �D�(֨Փ����Pq��Tѥ�τ��'`b��nq��c�7��v�#�nS��\V���y��gᇜCqn�0>6���yR%��=Qq����;���b#H6�Nk'~*ZNKITwE]6�P�-NB��L#��2��:8�k���U�&J�����!㭕$0��"Û��Z-K�=B�=7�8�R��M��G�4����>�U� *1>��H)Xt![ߠ�h���{qf�i8fg�b@�<����N���$���xc.�`7�zOb��^1�� 1���{�ZlM��,ev�%�HN�=���'�J���4�W��8�h/�D7evg�
g��*�:[V��e�<y�7/����`�m�`�P���i"�o�lh�n����b�+��.&�� (y[d��>�:����=�=��unP
�z9[����蔫�k�@c�	\��b6�j�2j�f��0�ve�Y|
(���A�	~:,ܜÏu���y�G>�;!Yy]&VaU�`o~v/����шl ���A�?�i�2ht�9'�4a���v�����n4M����с��Px`:�kd�h�o�v��졧/o�
Z�f{y��?��"��޻��Y~{���R��<c��zhj��|n�x�4<�Dw�o�H�~=���	�iև���~t�l���56ĉ��;,7�),2cw.��b�7ʜ���=X�Ř�l-t(���~��r��/��9�:R�4�����4:�2�V�_q}�l/��)v<�_żP ��xd�R��p.m�1�}qC���7���*�|������xi��r{I! s���8��	q ֌����-%�֟Fx�-%�˩����5ϥS�	/��Ȭ�-�����K�H��ܔ,��M�42���!�V�!l���YX� ���ƾ��B�W���|)�?-�	�8�?-��M���L��u�^�-rh��ŷ��2�nY�`ҏf�>�;V*9��	��ܤ�f�ۢ]���
�a��il;���������c1*����{��W.^E	4/1#XB\�kZ��^�+�.˘����ݬޗ6TN��w�[�)��j����>�C�9#K�)�� V�?�b� H�X���(�1
lK��.-����ԙ���]����W�;�*��qJ</�d�g�,��(f�ջ	�Aq\v��5��S£��\�6�����}��\y�޵�@+@T��a6�aV7��<�8���>r�9z���ԄQ�����R����5�u^��s=�k���N��e��f8OQx��)��x���u���?F�zk�n���0�Q	wn���`���_!!	�7	�h���_�R!q�Y��Cb�P�܇���6���}
H�Q̾9"���ඹrn�A����Y�s��+3�;u�Q�p4��b��@��ʔ���!B���I;�9��$!Uo�~�+��� �҉�Db�Ihf�=m�9\�E3IV��U�܌��mW�J	��C��|����Ԑ߲O q��4o���;k�^PM���I���E!��<Q(@i�Ń�+*Ɉ�<��-��qFd9��s�����v�YX_X�(}l?�e@As�:S������^H$���c���SB"�\q�3��F��ƒ��'*�x��k%�� \ �aV;2~�G)I��=i�fS�:�ŕ��@6�����
��gU�`䇈	�x��'Crr71S:n^A�u�8���%��!\����<I�����Ol#��3-%�Rv����=B����Zz�ũ�G%�BQ��_S�u ���(Lw.Y�8'H��*����!�ȐD��t�j;9D��m�NV�c��b�$��J8���..:`��$�F�d�x�Vn��� 'U|�ouqOg?P3vn"�4��Ԡ�Sƫ��*�$�c�x����ߔ  uC��wa�(L���$��[= �{��k��AVq��߿�hR8� ��;����޲~aD�����#UW�� ���f8����
�����/>C+P+��D���o��6<@6�`Qg�kP� ���O�ԗuE<,��k��{V�z|mv�1��T��Dr&C�0r)��R��[�)��&�6�DJ�}����#�,>�G>�x?�Lv�و`�Z��Τn���@u"1�A	��gv�N�}��A�x
A5E�,w�
5J!Qz�̳���̉��`,�F1t��<ӌa�/;��n��dʖn✳ǖ���Ѿ�o?RF�`\r2θ�ᬘ^/��s�m���d�������"��ڑ�.e��@�B�l�����$�$d2���&Ogh�+P�V���}�� �SQy)���E�)F@�@��,���!�U7�Q@ I�Bl�b��#Y(qP��x0Y�4d+R��C��5S���>3�����Ż�nZ[vU��s�t����})Z�CXfMU~ߝ!�bLȉV�2�r\�ON\�]%5x�R�������	c�?(!X��A�qS�ω	,�H�q#�S�_R��Ӷ��0cm ���!9+1k���n�����'
.
�>�*��m]�L�I��6���lc�bI�g���ԟ�}��.���m�	���n)�e/�<F�/v(�#�$���C�-e\���(�����,&_W���e}s�g����%
_���e��{tZ�"\�FBr�]wmr�}c�k�uh�'�O���z�
OSyd�j � �Ҙ�1�&[k�PI�Ԍ�P��D�a%��7ɋ�����w�3�^z�z~2�����d	�����r��^�F9�N�A�c�za�Db�Hsү��5 �0�Ɲs;!�� ���yg����aR���~B��+�T��]<ķV6*��Z����s�sd����;+Q�ƺ2���u�R�/���U��b�<��fY�[��Є+𞓌����y�m"��]�Χ̬h��WY�@�O	��ڕ0v�`߶ya�C6~��`l#�6�6��ݐ\."��k�~����`G�&���z��=���\����q ;��qߖu$}�/���b���귪Fn�L�����d}�j��0ڐ��r�8�9ٷJO^�ԕ�ӗ�ӱz���e�4|����������ѩ��7�P[\J����G�@]����?�<�uX�kƵ@��P��s�.ȪQX*��ct�[�_�׮���#����2��5�d��Y	 �� $���M�[ʫ��X��-<�[?�iu!��[�cۼS�>w�w��Q���T�o��~i�/x����1!(�K�)�0�CYDu«��˥��%�jfM����#�81q�Τ��7���o�V�E������F�00�͂�wD)�kQfG�{���4���JX4��� a�#A����g��2P�8w����N-oa|�&���O,��`=�(`³b̕��'L��hu��
H�M$�ڇ7k�4|��?�f�f�u&k͡������.P0���?�,K� C�`�m.��$�^�N�d�;[QH�ߵ�ٻMՋ�L��6M��?S��x�������D_v	��O+�m������ �_/K� ��Rݛ�l�'��߫�F�x�<�*^��o�o����l<&)nTw�ҁ��Ϗ�Rd��'$>5�Iӄ��^/Ϙ�!��)	r-%`D���d'�["x���V��8IE*��tR�6#t�;|��c)�xi�S���ne�ܒ`i�r�>;TS�Ie�e�-�&�Q1E�I�Q{��+D(S� m���+\ .Tg@7t�04����n�L���'��w�;s��d���jG�!Z��f����n�&������Y�]���m-/-d��e��٣��;,N#���o՘��8���s�MV���}���E��g����_��h�m/��!�#8�8\g�O���(��͂�꼉]o��*������*	CV4n�2X�a�P.�|6��Fŀ��I�#+��+��уwQo7����
D5�j��� Ą�dR��f�Ҷ����I�>*/�q�\<���
�����`�E�p���{V�O`Y�jNZv�.�g4��?f>�� ㍲T>ދh����O<w^�d�*�ש��	��<; ���{|
�Sq�SV�0�J�N���q���m(�;}8�6I�a���5 E��4Y4W�=���6���s453�-�<�;g��^�v�O�T�6�_ƑG,u¯����B��$$��,T�����R��QY��?)��S�QF�A4�����Q�Ŋ��Z��XF�E�mqŜ-��ְv�h��R| �XA���k���,�� �e��.��ܗI���(�[ �ւ�v���[��t��@Q��Q`54��@�c�Q��1���[��|�>]�m�V��[.-O>b�(ɠ�+(��N��aQ�;1��c�M��!w�M�}n���2]81�}H��'�U����[^}^*�s�Kb��H�z���HC4��y滹"d���WS�X=%.���%��� ��� <=VK��ډ��m��O-��:���h��� S_,�FB~��C5�<'
�D�H����p8�X���� n�\�h&�Y�]XqM,��i��?�]�硆u�����7��rJ�Q�*��/�ꟓ���a^���Z@ϒ��N���:�1cz�
���]��NY��	�Ã�<l��)Gg�Bf�y+�R��{�I�ǉ�FF�t�B�/�9�rFGq�lٲ^Y�bB�.ʖ��Y�ܗ�+�=�2H�`��;F��:�6����k:�>k��ݰ��1zd@����S�����b�+���	h`�Ub!`�D|k�*�7�$�m�d4��f�ފ���Ń8[c��o0�XM�ϓ��c�c���ʣ{�N����c_�f �c�9Lt�)(�/��Tk/�t�-8U�V]).v
��W��?��������`��eIdX�D����Gկ�~`�z��ē�M�ǘ�t��ݭ���&*|N��m�L���ĝ�a�xӮ�1XU���G���[q<SV��Iz&�S �=5{��!��o��b��/��b�T^��aY�fX^ ��xD�53x>����x�٨@��;G�9�8m-#\rx/8����X�Uh�w�Z���C��ϋ�n�?�֤~���(Q��Q��N�߀�;�,���w��\�3	�9�^�*<�k4���)��s��y�����')$'!�D��>���Cx��}��^0���z U{O���s�,�.���t
��8Fgm�/t
0�����t񉁚M�+��jAg�ZL��1D��ӞW���]��>'�(�L��=��k�s��-eR�厈����.<Y(��0�sIj�����8-��n\r�ʃ�i�u}�	�F�uq���w��@�{GM�0�	��/��*�;�	�lP�g�M�4Ȍ���J"E���J3*<�?� �%����#l�23{D�;QJ���m������Ȓ�Q����^c�n�,�%�5�3&A��Q�K��9��qީ@/ P'f����)��|��p{�1,
{��,o��6Qz��tU��u���u����+���Ac��9�� ����kA�j�{�'�$_h���M�Y��H�s��p^�wf8r�	��h�sDʕz��ޠjgx���-��̸Ƿџ{��Π�V�$�8�meu��윆���x�Odm���6o� �a�8H_*�
r�ύ3-q���׀���z
��Nc�u?���P瑼�yj�|��E<��Q����$����.����\��R��a�!�z<��Qk�͆�=z54w�p:e-9/�<�*?؜/�4��	Xt�|j`�9	m�w��,0@;L�[H�M�H�h�����;��/����e�3�~Q�c�`i�[�C���I��1�d؉�1�}�2.���	_����FO��K�	���f@��{MD�V��ή6Rx�G�RϹ�������H��_}��t�����{�_L�<��}�$�� v�iG��EB���c�h`��};.K�� .ڪt�^cC+�y�k YՂJL� WE�D��]w����<;�jዯ���Z��^ZhP�����Њ>���Fƌ8���u����r���1
e����|��*��@Úx��_��c#H�-(uf��PԝY�EU1�.<�%疞sŸ�-�N��Z_��ӿ���$\�g����Tv?!�8��d[��=��]�\ڢS��w(�I��q^;w/���,�f�����;C��Hh3�%��ԇD%D:VX}�_`�諢��½r�3����}�=��H�ۛ���!�ݪ�)�����e� ��A�&Doq;�r3E�O�ݦ��j%�P񅹄�s�� ����fkSY>!�ȴ�aQ�˂�[]��ڵc�� J�H�ک0�_�)���mZR�E��
�'�頃��# �y6��in��9��m	R��yq�)D�� J=�lf�5��ِaz�ٴ�},l0E���벩�����G,���I���ů"b����\ �u`l��./��aT��(F3	���`^i�,.uK�B�@o�})��!W/�2R���z����T �C��o�⸃��ɟ���h��ķ1V
9y�#(��T���Q��3��NE�R3m�!���]g�I�����Ε�{xh�w�7$��K��$�I^�$�� �Fd��v�d�0�J�AQٸzX��V���}#�d{q��و��;o�(�y,���}�l�����}�:�I��G�{: ��ˮ��[����w
_ �a�3н���FF�CW[�D���J!��Ȋ+�Ye���@-�%҇��:D���Q��9o��J��(T�@Ύ��Mo�*��B�����������R��GV�p�������G(�O�4�-��x���[��U^h?1�R%K���x��?�R����?Goo��+��c�B����T�x��xKV�r&M��ѥu�?cI|��U'�I�2)��nA��t{]�@m|Q�ӹl[�Q�Q�ܢ>�lL^n�a�פ�:��O�Z*�\��8����1��_��w�74���s���~t	`�	���̋c{�ȱ�j�Q��-��љ���H���r5tƑ��f$0'��u����7����4T�#4z�
��{���LSX����O�s]gWV-`�����PtE���ഀ�g*ݟⰈB��|:����������G�1<���Y�W���SV��Z�u��!��S̠�; 8�/���b��/l�����[��RǺ�ׁZ�<5�r+��v?¦���c����>+�|�lN�Ë��M�SB
ZJǠ�4��):��M�\p��~5k#Fd�#�3���z�<$\��f��p;���fjܒky&�ƨ�L\")�d;C�,����F�^�B4�B:ŷ�(�0�^���Z\�.�(��������d�~;J�ҫ;�F���gjM:�P���K��5XK���������) n��7��&��9[yn�����^�gG�(���X� 2�1��L ,d�`�j5B�<^}>D���+/@e��M��k~mu9�ۇ�Mu7q�r�G�����@>NMf����>	��p��� +�*�/���]������bq�s�s��E��tz�Y%�jR����0-R�4
���^=��22�B⩶U��y$���Vu0��éjT�,�0���p�,�y�)1��2��c�i��ŮK\@D����P&��!Bd�S�`��x#�`pzσ��7U��� �ފ��۝N�˗u&� ��& �I�tV?/���fZ��&1�<ظ�`��0P�@#T�":��1ܫ���嬾z��9mt���|��]��4b�ƙ�*�wK���I˯�	y�f��Ϙe{W	�;1�_�����v��꘯n�/��y@�b��Ib���`���˟���*��@L��)�[���isC��)g�x�A̘�G��v&� `�펕�8rpߪ�\Js�n��->M�&�� `0x��������N�*����0�ɤ�V]���uh�ж�]Y�&U�!�p����9�"�z`۔jG���DF��,���EO���d%�H�}��`�c�գS" ���С�Fd�>)r;f_as{qW�C��*�8� �7�}O����x�*<Oڍ�/�α-eWl>�eyr-��fuI3���� E�1�p�);��J�%Eʐ�V~��P��`�Wn+�� ���vW�����5����ܶ�ro�y������I1o�~�(�p�Z�7uA�yUy�X��'Z}G�zX���m��?�~����`���V��j���
4�|bY�Y�|y����5Jny���X���k�o�'���i.��8So'�SM�}H�ZX��y���|��1D�H\f#G6�V��1�7�}�ۑCC�n
M�)O)���O���o����P3s�YQ�,yM�G��*�,��H�+Ա�n�/Ɂ��E��M̔;�����;~H��v�^ærm�ӖiPߙ#�g��T=��'^��d<h+�,^����V�� ��S�!V<�a0���;�s%I2�#ٚ��k�� `C�pY�\��B�C�>��j�D��v��o��I���ͥ4�Q�r�u�Q��d�n�ڕH4�Bt��QSnw	��ä�ț:cI`��޽p�{�����)�-u��>�㸅��5��p�&�V��Ä
8p�	���Z����,�z�p����֘�)�!�Mʎ ��%�5@�*t�IZU��T���z���q.T��i�Z@�q�}�ɤT=������|����X+���i�T�^]�,h6���D�C�M�yB~y(��8�_����"��={Gر�^RA��t�9[#�J��Z-�j��1�'��w�����1��n��u����*���%�8V��y �V-P��
h�;%�kl"�+	�$@����Z�Chf,i��#;�4z�^I=��J�X�u%v�ܠ��B@�%��jD��!M���&�X3s���F��\�#a��"N��K�Ft���j�vvC~����6�x?{0V����?3���d�dh�J��>��qln���q��h�!�:En�5��46vĝ �{
�m%�]����Ӧo�E7�.� �s~T^Kt�EDr�6��o!~G(��J�h���[L�w���X��٢��8�HDE�컾9�ϸ'V�B�.��թh^Ȼ�%Tp��߶��Co#�(��S��>��La��<��	��Fz��A>w�ع��&��$���{_ut��/H|�}j�]W_����ܑ�i�1=��.P0J���9���.o�F?�[��fnD�.��>�+�����b�f�	1Ail�RW7�>}�-���vsb5ۚV�ل��p���1h=�h��ܰ-�5[�,��R�9>s/\΅�O���T-㊁�?��v�\�	0�'\��z���@t�h&�f;�@�*�/rTo�M8*��4�<!�1@��؄EcYu�����1�-���>� $;���t�8(Q>���	��)���i�&޹���Z���l���^mE�k.
��Y7�>�n)RE����S
��d!ȏ�"���q׽ͭA��������>���v*V:��O����a�f�8:���f�{9��Ӿ�)�ǹE�_�Ԓ���U�+j��K�&]���H��N
���M�����]�̀!��7-���Xl�N�f��:=m61�_��y=V��=��<�7[�SA���b�`�r����	�=�;�-
��*T`Ws9j�8PH���x��TO]x�N����<gӅ#P5�,�ό3 �l����]�����MC��4�u��Z�^�&F���P�f'��j�'��ׯy{3n�]�v��*���љ���E>��.QX^���F{� 1�2YH^D"@�'��v�>7��&�?�N�?J_X�=ei�S�ms�t���2F*V��c���������2|�W~�A����Sx�>�	~��2rR��3b�S��f�������+�"��2c-��{t�&X[����&�0�F��#����֧D��6T7��--=�uO��]�t���f}�z������u�F������2�[���W�E�ssf�k�!�
��)�GD]鶟��� R=�&�HG�j�l>P�瓐�[��
�mt��^s��]���D>�дh���X{�
�/;7̀+}&������2�2+���[yR���\V��#���Z��Y0�a_@�[�\|pȏ���c��W���?*���"��-�����$dS��'��K'���#]��:���v����`���M��e�8|Qx��T�K	��W;}��}6zǞ	O�q/ѽ$C���0"���>�%�O�:���V�?�� 0b�u�y1�@5�)�T��f�����_3B;��-����#�y7#m>zǜ��� ��B{�r�^�����Ж��SB�-Ex�o6B����?\�$t�K#�i@�#��"�	C:����<�z5������m
����S|}��=L|bI~V��Yͥ����I�.2�Űv{�错a	�R�b/�F��
�!�O��Ԯ��&�r��Hմe�Y{�֟ñ��M�������"5װu�?�s�p�[����B 9�f	t?�r��*c��U�L<��2P�LH`�}��>��|X�3H����A?B�9���y���e����L�� �љ���^L����0l���v�)7��$9�����(T��Ŗ?>ZՅ���X��P�����l� J�恆[\�y�E,,K���=��o�sų!��Ŋ�⓵�C�t)j�fј`�%c�[�"�N��Gu����̗�s)q=E/�T�ﮛ�*��;;˩�|���B���&��P�=����(Z�"ȟ빿#=t%��r�IK�I�Z����*�O*�;�;���Ӈ|n�ȴ;0��ī�{q�4. ձ}�o]
�:Ĳ�kM?iN��@��iV���߽��RZxVE�i�̋�S.t��=��A������k�K�cYY��fU�U>�ߢ�)-�f�f ����F�ɩ2�:�9��6(t�Ot�߇c�E��%�V�;���l<�={$O��gB�G����'�1���wW�^����H���잼���	\�҈F�ù;fĻmޝ+��������S��D��cK��ߺ!65@Ԋh����,/�B��k	k:y<J,Fs�vU�2Q��l��x���-Iꁍ'�41");�8�&��P�Ix�Q����EI���/%{7�\A��׷�,�C8�5;�-"�� ��P!�]����6�`�Ϻ��x��*+H�ܫ�kn���Iu8(���o��T�;LKAj@}Y�/̗S�8�p]��p�S��o�A<l2���Q��ܡ	����f�t�>P�i�+|qR?�k�F-R���tu+�\w�2V���������L(���H�A�)r�
���(��	�-k�����C��3%9�UA�M�W#�P�{�7�X0jGf ��&"M/ �Fz]��,��.�(�.h��O�Ѯ6���,�����\/W+���:8���]��j����"s�o�b�EK�M������BN̵���!Q^�-G��T���NY��ЍU"-.OZ�(����tCF�9������z�-�z@����*_��Y��տX��0QI�l|�g�sҋ?�=����^���c��f�H�js����.Q�"ە�D6)��]r��V�G-�e��_B"%8UcA-@���2!Î�cT���^}��_UM&kV�M@p ��*D���P�b���p�kǖߺgi38�k�Y�ƪ�����>R:U����O�k �1f蠇��n���\au��/�uH�<���̙F&��~�)���
��#�?{ �l@<�A�@D�Z|��K]�@��D�� ��1�n�s����f���bw��icX8b�y�tM���f����=U�G"�υT7���?HN��E���c�{�r�ɱ�G����1��߳������7ɃO�����7��8�����!�=�[�X��D���4R�Zѩ'��:-�4�n�+J���k#k� ��ю��Ƅ^��N��V���_�|�EOĥY�_��n󧕾�Rl��4�s,@��o_;��RO�y)��x�_m-�7\շ�+wt�ɖ����YX�ݯ���9OR�/��3��5��9�˦+�-L��"����ر���&6��4!+�I ��X�=v� ����J1E�I��Q�i�r^��i9oe=�f�3��I�zi�0L)���1D�}����f��/��u"]m��M��w4���{n��vG?�X.T\F3W��y0ky��!���":�L>i�ΞBv��=��8��((R���*O#}�-�p8�z������X�I�5�A�>���ETQ��e�Vq-f5V7�Ep�=���X��9f9�\R>Ĩ��H��ڰ�D��p�)�PՃ�Í�V��)�m̏_��X�h�c��K�\Z���P�ޕA������u:����̽l�D멝Fτ���4�����x���g���5���)o�ٰ��@�2��) ���܀�(���7ƅb���Kb~⎫�Kv�h�(]�;5�?0�־�)��O�����s3��zπk.�F�7E�j	;��`�6��Rh7�Vp��O���jT&���eJ��?N���ā���v�P�z��G\�#�1�М�e7Ȏ��v��"Txܾ֠Ӷ!��J$gH��pR�sh���<��-�(�e��c�vZ8�y;��}����K*8��(5ۀ[�WU%6^���y��?Jw��?h��1�����(s�9� �9qL� a C�۱>zd.�+��Z3�4�Q�)�Y1 +�7;�3�b�lۙ!s�]�ȢXw9{,����kR���@z&��~6��^:�9�?�y��\�S�j��m���[��nh�׭*��.�v��?��\$�S(3�!OG����8��VeC��;-�K�`t�:wig���J&��C�8a���Pܫ�`�/hpsMGׯ���N�����KZFl���b%EVi`��pBP̰E�i c�J#F��K��A�xL��S�#/ʼ��/�Z��e���QN�0�ڕ<1WIL������;d�=��grn�o��εO�V�����+�:�[Fo����Lݷ�q��dC�渉eQ;�qk�pX�8j�Ҵ�!���`��y#��:�U�ʲ=�@_.�8��zXg^\�M*�� ��6�Q3&�����U���6/|HUa�H�q RJ]ƹh> ���B���~���'wÕ/��?C7u8;V�\%�&�"���Z]e5�&��_��,6!�S��;��qi�q�����"�C����a�]�2����r�/5����*�\�����37������FէE�����2�(3{C�������l�s���\�m{��'E�/�U8&�2��Sm���Ʋ��K�O�;%�.�гH�V�g�����K�޺LB�2�Ŷ˂V�u�]*��3wQjƲ��=�9g)�����?���,sG_� gM����U깦��.�	��	�(��[���4$.�9�<ɾ�L1/Ɛ���9��>�$�`�Fn^��)[�@f!���p8מ>ۼpMjY tqFO����T	D�=`!�Zs���_�!��7$X2?�H��(��r�w9��2'\V�>4�v�2q6��R���rD��-j���0'�D�>;�.%�5����h�8���n8�sRu�����N2D�IA�u�Ճ��g幡�
B��� �5^`G�-P`��Ч�� ��=t�Q^�a��R�kͥ7x�(Ϫ�ߔaz�B�AD������⮯�8�l�1��&N���0i(D_eh椝�o��zIVF�;j�i����jT�?���w$5��R�d�s�d����1�ڛ=t1�Np7N5�T�5��$ת�(I���z�(g�mV�6 ���h^��K~e�g�DbLc�*RdM�f�M���*IY�������w~���ۉ`{��&�9;�;A���|7���~0�����	>9FdD ҟ;N�]�O4�Y�*�7�,{�%������f�rb
D�P�K�c��{qǊC�&[�4L89CĄ�j��f��#��;Q>� ��j.[��G�Սͮ�=�Y_�g�?���G���c�� �&MCAEP�Ixɾg���/VW'��F�]ضL��y$�32za.�z�T{�\�o7n*����:��������˄���E�4���E���昶�t|A�=��X�ܔX�:d�|y���Ë>�$@݉�j��zCr�
�%-{�:7w���jcu�?�W��*��~��ŝ���ϸڀaw77I����C�_���u��Ev�~D�v�w�,5��?�U��/*�-7Rp�ʹ��b��-�3�v�Ä �K57���u�����J��F��"�5����]ٳOr/~�Ns7K	;�O�E�G&��q{B�y��ؒV��(�r����
3�e�J�)(�ń��`�oJ=�[<`Q�F%g��J��UU��w�N�-:���B),1)}[,	.O����c�.��p	ƉH���Kp�� ��xtqt'l_-rv�՝�Ɔz��ێ�i8�߾)s�E�-�&�eV�H�j�����^]�i0�m��W��6��!�<N��uGC�ٍp�7��M�AG�_�DՀK��[ @�V��X��8jN�;(���'�ƌ���Wk�O�Yu�R�,n��9�s�@�����8���֬
�@�n��WU�с�J���0Qv|��kXp`6�U���&�
w����_8n�bˠP��1������\��p�-Y��{Ĉ�)� 04Ӛ?�_=N�+N��,b4��+�Q!��6�|��q�c�xW4�̟��{S�L(�!�%_�%��$�X�Š�������j�3Y���D\f!��m��R��9\��:��ܤ?�DR�u;��(���걑��\B���h|7N��
���`ق4�^K�
��R�5Y�&2��.�P6Gqw�J}H��/���Ј\*.[�~`��R�q�C����*�v]�oW΂b��yM���b�re"uܑx"������Ô��K�;fl�ڧ�h��%%��u���+�*%���j"�tqa�ȃ=5���&j�w%�$�Q��=�L� 6��>�ޒ'vq�4����B5��/��h�bI����+/�I�WX-�C�i{�<���#�w3Ϯ����H�@o��cL�Qz����-��&�B�9-�˔�In�P��L8.�.�$����yD;%5���'}ʺ�`�T3�������b�0Z�##�����#]t{�X����3%>���56&_U�%s7���+>4��ϠlzH���P�/�􍿾�b�ⴰ� S���wU������U�NƱ*umR`ؕҕӻȢ֚gY(�Y�C�2	jh���9�Q/w���IX�r�є�hH�y&�{�BR�{�����/�a������BQ�C&]�]�VE�����<�+b�ʑk3V�x�"�/fԾ�{�`����b�����k���K_��kqz
+={/�� �c7,����Mm	e�?E�v⏦����ׅlҟ1C���l%�
�Wt๴��SFi0b�4�yn&|<�^��:>�O��=S��H/L��K����/Z���������L���r���,�L�(D�ʻ_��LMo�_�\���fW�����a5��S�H);�xCBPG�]`�ϙ����q�J��V�8smp�D�0�����2d���^���?X��jz�)���#sX���d�t,��6�W~����y�wv���_?@XA@P����%�r�Ux��F�J<u/�=���IG�㸶��lUǋ���c�����HN%.77�1���T�I���l�FI^\�XTX4!��W���.UpY%f��9*t����]�T��-�/>2q��,5�_/�����!Q	C�!���7�"�Г��=�
S1�3��|�+��S�ki�
l��4�sž��k9/��W+�ri7�E�+7*vw>�r1���z9��}�-b6%�=n�"pJm���0�8���� �C�+��'19Q�E2�ҷќCu��T��^D�~�s?[`�/Ye�$���n֊�O�:�-\��G�vo�Aɾ8�hv�پBi��� 0z��'�A'�^���_�6 Ó�~A"T��n̰M>�<���GL��n`��2�Q1���D�D8Y��漍̤όZ�h(m�)i.��#MrUy����s�쨍#��5|�4��ߏ��7���7UR`���֏�����F���f�����G���4���p��4h_8���Q�>�]i�3���e��S��o�e#��Tr�.tAG�>)d�����$���v_��!>Ps#jڇ�����+ET�m�g
�hzY`��)|�T{�4E΄�g?lE�o8"��2 s�C�Kʎ�ȕg�Ȁ��H�0����uG?���吻�����MH;[O�z�4���v7�5�x{⏩�$;�������j�`G�t���b��S�b`,��B×%q5С$��Lq�M��~�kʬ�,�<�P�ſNC�%+�N7���D�en��6p�4�^��s���)m��0d��z*�Xö�Z��UX�u�|*�RP���D�F(�3�����}O[Ml�P�FY����_9���� �FpI�2�+L�@K�&��a��6.�7g�����dڍ_�Q�ˎP�S�M��3[%��>�����Fm6K�G�ǔܭ�ʥ����ɰ�m�hӍ1�����I ߃	ެW�u�/�I����!8�&��j�5!�:�{�Sj�{tIx���%[Y��QE���G�I�NJ�Ղ�4���)�k ���Å�����~(^P�&f�FTf^w���h灃4�2U)Q�l���f�|���B��AiA�M��f�j���U�|�0m$��p6ڒ���8�v�M�4n����*�}]z!�IgD�U՟��@<�8��rY�����٨�s��?�	�H&g�ޭ��F�S.�<a��+隆]�� �93�i�	G�2>���$�I�������٬�[a����DUQfGZ�6���s�ܐ��W��܆�A�L��0�6Z%��1.�H�7�(n_s�� ����z�8�k��"�I��d�f�8�C^��A|yh�Q4���ӿ���q�G�"Y�)�� ���L+߅��SAk�]�h�h����3=�k�.��i/�i��*@w/�n~˃I�Bn��8��6j�l�D@�Gs#�iC���~	gD���c��:��`e�\h´��Lք�.��zl]�{�B�_���U�%}fS@�����y�k���SoT7n��.w��̝M�T��o�Jl[�(-�9�8�@J�p�ɏ&�sw�'����p���2#3f4�u��Bz���r�;N��ͫOD��n�mtc������ٻ;H�_3c�^hg?_�o=�
K��;'t��~d8�~�M|xǻ:Ø�z[÷�f�oa�"����X;u�DO��-���H2� �8�& Ң�W�c.݄G���A��s���IH=%F�jd3�3=���o�����&����WFpv��]�.и��4���(�6���M5+�������]�yu�Ƅ^`ष��+Y�5�Y�W|O�����=�aХ�� ��4�����`��w�F$����2P��ݣ���"�� �[AȎ��ZL|y�ݟ�r1Z7l��/�qX��W
5����?�/ve#�W�*2xޞ��;
�9������hZȜ_,��.I%�D�WVE�ѳ l�������.�r�ü�����[��u�(�ķ.��vԾ�>�<��|Ѐ-�E�\i=�cX�w&'��>��-�p�����y��Cp4%��Q.�k�ͼ}��������`и:�}R�n���A���g�{��i!���o9���?�g���]>?A��[��1~nޥ����m.2����z��lٿ��y����} !��[�o&U�Sv-�V귫,9�ک'f�y����5���V�}�(�3��,����C����E�6}a3хar�A��  �����ȃ��#z�Q����M��'� SVMӍ������
2��.M�\������l��*�?�
Gu��ʡ�4K�.s�u�J�D�Q��I�wFD֒�Ɋ��^mZ�t�W�[3��7f}�����p�c}�3��)vp��u�a�	@9���h�Yh)^c�]v�(�?](��l������H��[�����%�f�I3:0���N��-Ws�ļ�pzS�z�;��i�F���Ji�k�4��s�&�!����V�EᎧ��W�;A����g��恁�wl��8�|l���6-v�����fy���9&�hl�*&G:�#��D����8�a�؊�7�)�����6�b��v$���e#�GJ*P�Bh�W�� �w~��9�?��Bz-Cos�N��gVY�|�1W^f�XȩX#��2r�pZ�&1Q���f����#��p��e��D�uȏ�1��� 2rm=��@�U
��ml�0|^��5�r���T��TuҾ=}/i��Im��,H���LW�S1{<D�m\tމG�;�+ξV3X�o�ͽ�V�=Ǉ�AY�	=RyS(��E����4�A���&Bk��̙51U�࿄�8���]�yK���8~t��Z#uѰE4�������x��x�ٝ���^�x�o����b@��9FEď���I��ܦ��
W�(Ն��(���4�7A`Yd^V�Qo��#��,�mR�Y8��� ��j�>R���;)��B���q1�Թ֟d&H�SM6�+)2�Z6[�G7I�Ůr���p|�6-����U��M�
�!���k#�֬�?��)Ϯ����'D��[~Z���FQR�/�����e���vL���u�!���e?%«��\N_�ݫg����S3K��kf=cZ�V#,�m��������b�T�P"���N,V4nq�>ϙ2�ΖO�5�3�_��x1s��(����k�Y�9��mS����,	��K�������b����̧T�_��� �8^:tU\��̠�Vg$�
��Y��Ȓ)�<:.��aho�d ���Qe����ɮt�-���?�&�1㔛����=ȈfMX�0ݘ��)\���4��|6E��� �a��T�G9 �����@�!�%b�}�)&2�*�P�fX��f2�����u�k�Q҅��Z�H��S�9�|���&�8|��#p����4QD�#ەS�,���>�a��q��x6&��r����':X
����ŵ��-�u02/��3Ĩܝ�o�x=�TQ���g�l���q�:��E��������p���@�$��{ؔ����8gO�AO�D��+�z�VCڑqj����3Ȩhu�j��L�I��߆�2��(q�o�;k���cZ�# 4�xˀU�Km}lZ�8�u�����.;`9�]��,�l��B�f��,�%�ʸ؎ԟ<�Qu'������'�IV���ʹ7x�3���$F��1�+%�*�Yk��L,���8�i^��vn�\�{�{��Q�7��h�̠��q��K.̏����6B���+Ib�=X�s�VA\�`(㪜U����{�=�3�uf�{C+���U�t���L숶+�#ĩ���r�3�yc`���
EB	��.5��b0jMl� ��d��@�]��蔲}�5��h;@�e*qG�	d0�|8hЌ��!2{^�t |�1����2�	p@q����R�T�o��6y��&��*�E��8jф��u/�Ŷ��~ہ�I���}x��<�����A������+;���11��f_�V9�;h���N�u�0[���|�����W"��]��ڄ�[�n(
�T���>�/��o}Zt�׹��f���k�g���&|_�X̔Y�E(�<.̵-{?s �B�iV����A��GՅ�� �_�l�ώ.&��� %��V���0=�o�[�ڗ�1��oq���<P���t��`��\x��W0.���=!�_����J�'p�Ɉ[x�u���d��2�Z�<O�KtbS�8���?���O����Q���uT\dL��Bzl�4��E3�������T� �1e�.��N$�n�t�	�Q7A�j�ČT�j܄q��,cхj�z���A�W��FN��,JOg�N�Z�b��&l��a��1 ��"�#��ĳLؾ��a�w�k��~�")�w5r7�ښ0

�H�go$�+T��xqmQ����u�7�fȠ�� ��� [�W�j�љ�ː�YT&�׊Ie������9��B��W�� ���k�;?ҫ��BY�0n����4�ˀ�����ֹ�"����b�g&&<z?�a�Y�e�*/��^M��y��m���D�-. �
��7��� �-~c"�/l��FHע�'��2��R:�Y�����O���*�7��M�©��n�nJ�]�
��w
��>5��C�9+mٱe����|�#?�)�@�`'�BxX}}5_��L�yo��������=d~�
��=�!��յ����?�"+��u�h��%�^����'Mk� �Z�M�N:I'����m��߃3����n�n+�'p��3��2P�%#r���.!���9�~
\�|�<&@��!~��6��d�-x�3%��lʟ����X�́��)�g�Ll� �t�I�#Zpf�sm�Z�����o��q��
���u8>��C��@��g����	(h�:�T}d��w"����%�w���� �&_�K`��f�k�t`��o�����k"@��0���0T��X G6�Jy�"��B�������W��*owQ&u�g���*�j��鴵������0�@(�A����K��%�`N�$x� Zdf��M{D��J"��:�<qmmwK�����;sa/+?��BY�7j�E��*���a�-Ɩh�zҾfRs�v����C�Hvbt�=l�)6r���e���rU(�t��V��R�}��C�B;O硯�Rg�4�".��&U0���]�#W{����O�ݽ�7�^Y#PM�F��%����;ͻO��e4���iFxcr�-r�;#�cy�~1UUJ�*Ě#��~>���,��w�z*\��/z^��f�&r��޿�h8�J:$��oӐ'6!�mu��ߘ�3Ϝ�
�2�Ci���
柠A�-�)[��=�o�eD��i66�̹L�u�
g��~ 1�a�	,�(�RfN�Φ&k���吽�+dx�uT^�}7V�~��WEED<�wH��8��18��?:K����j�I�P+(���z�F�Ҿ�蚫�9��խ���4��{H�g����s�;NK7�&/D@��fF�:2`q
8V�t:�=:e���5҄�oL�;�m9i�˕��NO]�B6��i�n��1��vE�k�.�JN�'��n	�uv8Puΐgm��T(�^�X�@Oim7�v�Hl4%���jel�M��5v��F�( ��8z�y���~��Be8��$L$-z�6yy�hoۛ^�������C�(/�<؉�Ȧ�shNƯA��tkGP�97��0b5��?����	W��@,�s�{MŴ`�u��	��h��¹����F�(�i�˰����j����c����󯺒�D� �~?�6m����]���W�W�?���}��ƈi,��<��[��փɃ����c$��)���Jv*�9wK֐�u�r��
3�Rbe��x���q�1GI�E����6�O�$�0�f���&��zbh�<���5�2=��BR�C��3Ȋߖ�~�p�0Y5��Z{3p��Q*�<S�Z��t��:��՝_"�	�pʧڐ�Da��1���q);�軇��6�1�џt�̈́�=�J�_�dH1��I'��5�"G���6{d�8�Z������\���w�M<��k/�����X`�P����Y
�:�!�8�m��f��]�������PTg�;?��W�QA'���;Q�4������?�E�|���+zl�g��o�s�1H����,[p��ˇ�#�t��n(�u�OY�v�Lc2�#�K��#�q�ã��e|�@9��%�A���buƠ]=YΖͅHt�NR�V#E��
6��%�	�>���ȁ6�eŦP�|/����3�Śv�Y�&��`w��5gS���<� �����T���T�-k�%�E�m����+ٓ����ͫ's����Sw���p������"<�7���f.D�R�7��x6�\����w�J|�1-��X�l�*�@8��W@|���_b�aS��㟣�8?��EW�2�^V��2�� Ű���C5Do�vu/Þ��a�l9���_~V��m*���c�Se��
+n�UbUܫ����%��wuMP���� ;ٲ}��"7o�<�/�e�N�?0�t��g�iЌ��	��	R|��W���+=��	���O��&ފ�����J���H��Tz�\��We3����u��C����pM�r�1n�����%�z`� �'�A�n���5Y�t�s��{H4���UB[��p����1�BN���ZŇ88Fi����:%tS�e oۧ�k��i3k3u"H�ҽS5���IN������Sc_�O�����+�ȩ���u;Eꖧ�u'��֝�B��$c�����SY�PnS֮�r���F����F�O�����(�&f�(�~���x�C]X���ݺ��f�N������'/����jd�!�bG���X/;�����"u�{����sZ�Ʃ5���֊9Кds5�ej2���<\��Q�v_P�� 0K�K�lpb�`]1�|O�3�u�-�/�+���M�w�%iO���>��{\����K����
Z�S�s�5�*����!�����|Ν9ϔ��q��
���&�'��dт}��N��sϪ�����2�O�	���ն>ڹ��| �!-7��}2tkr�L�|kN��/$�N4�>�̩R����tv^$~h�c�;4_�Ht{8�1{mkH�")�M-��*���I�ܓ�D"Q�9�$�x{Y��>�J����[�X�?���0�Ƨ����4x��-0l��|<�ʟ֌�GY$����p����J��s V�,��"˱yB�MŉH��p�w��=0�O�%�����%��O�j4a��fļ�[J���H�a��F��]��{�d:[e@f�o͸��S:'?��L�M7��bt�N�Ux�x�;�lb����d�R����3庿>j�a�W8��"��;���ᣇ�CQ��@�9�Z��)K#��Y�Oz�_��p�8��A<�!���g�+�B����=ָ��풃�X�҉�G�S&�2�;Ju
�ry��ol����Աʹ�����C<�f� Jz��Ξwt���[��c<�3�5&-p�4������5�鴙*����<�#�J��ܠ�
ƒBCЀ��[U����w��
�
�7�n�W�%')��u7ֿ���>��E�6��uN�M�	����1�P�]�c�i�!�y{T�ht�P. ���{I�&�Fy���!r3�E���Gt��Z�<�[u��P��&h�\���2jl�;����Ӷ=;�&�r�*
to[ﯕ1p��-U^B�+s�Mk��	?�o�:!l<W��+֒�/w8���V(�+������Һ�%G39i��c������⟆h!��݃4��[�}q��K�=���*8kJ�L���61��
FtIA��o��E��:������__mG�HT�����]���fy^��LF�H/1��z6�~��<y����G�yj��
$���NlʩP���e����.m�7Ś������hԢ��&�w:�-Q���*%b���+�#]���ѭ��<���1�m�lc����"�5�͙���x�egXQŮJXw�t�S�X�?ncX�x� ���/�A�e�����ȇ�%
;���%[��M�z����A=���Xg�'[��_�e�-w���/��&x�bX��&�����Q&=銩�c���a�,I��"����S p=\��$*���M�V��f�H���2���':��-��.��x�ۆ���$�����0g��dX/�0�3���L2'���J�A�����j|[�	��Ј��[xO���l�J�1��,�P'����G��wJhV���n3��cu*7W��]���u���
�OC�	�d�7�9��s�DvW*�u��f*Y���~�G����0�z���d���r'�t�r��k�ܳ�8�`f�Y|㸆�~7�%&5t���9�{�+~Į(��S�oA=?f�`�o'\�;�
�&�$Q�s�x0�������X�s����<uի�˞�4B����,g@�A�l��+���m��WN+J�F�]���5��4�-��?r�%K-`y�-ŕ�%H�G��S�)��n�ؖ�g��a=xt�4!����}�`ayV^�
�vUq�ét4^�x�q���'?PV�?0��\	�X�/`���d��bA�h��ʇg�}h�������AL�����e��c1+m͚%o��L�B�_7�2e~7o���E�o�����hc��7yZ@C�٭�6��([��ME#m��4��F�w����%9�'�{3�'�c�h��1��˰��1�[��~K��M���X�@�➏E����q�(�%�x�|n��)N��%&l��J�iCʨ�)p�F�{؂�a`�i��ը��t٤;�cYB�]ɴ<9uD��\02�Bt��2뾖*uH胛&��S���Y4����$愋�w|��ǘ [����P��+@�B!�����E4�s�F}��H����8��>�Dq��c �J�z���$^�"�^��k�$(Rƒ~~��X��;w��ɘ��d▭|WAR����x��ED�- ]"iE?��^���@��C�g��)�d�0�O_+Ǌ���p��U4�ך6\`I�h���7�����O@�����q��>j9+E�;9�O�~�oI��us'B�7թ�]Y��C�F�QiYJB���p��l���!k�hJCML�#Op|�D⠂���RX:�Dc���ix��z��a �Iٵ���8�fUiq�u���ƚ��O=T�FJEi�qf��U��xQ�W�1��""���`&���Fz�]ʆr��>酇[�3d�ݴ~R��Bڦ%����m�4��[���w"�[���� N��L��\If�~-#�ü1��5������r`��8�� :��-��{���8���4's�S�t핝��^�6|ɣ�:���<���q��?�t�/"�ـO��g%�M���E�?�rs�R/�wZw�����Y�a�Y��5�W���1N�@��<w��t�u�	����@��4�&D�ǲ(`�f]3�w}A>�ʐZH,p{4O˩)�XJK�c���i�����i�={���_�sے�)�˄��'��k�%s,7F"}���z�����f*�1��K ї�w�󃦙)R1	_._�m-Z���o�&ڻe��l� ��42u{[N���L�Ǟ-ʯ.	3�ꝯa��ҕ��љ����B2�׮�e�<��i��f�YTu�(���#���Z(�����`DA�rON5��#[ͤ�N�N6U;B�������v���vqԔ��a!<�\id5努�9B�i��&%���~�#�4���'���v$c�PO���*���"��
��R��80���7є�"�R-GP��f�jZ�)�R����;��R��(΋Jv�a~|<���Z냙@��]��SMz.���l����W�b��aoB�@����ldG�Q`�/u%BL����\#��پ\Į!��W�S���k���Mu��z.C�G�O
��yg�PHJ�}b��r�8����4b������Gf�{��Ч����W�Ta�o�޷%P���v����f�@ɮ���y�f�%_C��Xۨ�umBïJ�`7�M'������D�@�,U�������8� G�?��BLc�g���D(XN}:[Y���_����TUF2���m讛Tig�����D�kW�@uNC��\�1��A�a�ۃ����7s�>O������q�h��g>t[x2�P����Q���8א�H���_�,_����ކXq�u����R�<zR�\�]�$D��t��SHY�������� 	���mW'��Wn��Ж���2U�����n����M��V����}��;�c0�nxWA�����%q�|��Di�K�j�R=ҍjL,�@�b$T=�x�Z�J�����X���J�s����$R�����(���jc�q������O�o�h�^���`��U���l�� ��+m"���C�l�ai�L�V����(w3]$��"a��
OL����!�ޯNS�-`�N������ه`���� ClyI�8L�h�Ą�o�h=�0�O����b�jLk�k�M�C0�@�R��r��a�C�� ���q�!.����_!iy�k�p ������Y#�U�r��1/:B��������ӘR-pX�g���s^�s�����i��������Gz�����Z%<0����`��%'��Kd� �˸C���e���;"�\}=Oژ�j�㠝u������v�e�%���f���l"�����<��i���E)Q�E%������4g'/u �8�ch<%�ț2��͵C�=R�	@~f�o�|G��=K�p�B�<���OQ�o����N܍�é:>F����Of���G����^	-�O�\P�q��JO*�ϰωK�Ɖ�V,�� �0�<�`{tɑoW� �䵘��j��q���l�)�U�^������)s�P�́e% ii���Q��5�h�!�4N�{��cF��VY�4�y.�e@J"v���s�P2;s�~�,�4U�N\�'���l��ẋ����&�T���e;P�Z|p=z4�~���f�ŅL;�WѦ��vk7l铋(�P���a�-�!T[N��j���ch�
D�gL�.�\~�t�D���U��ѱ'\.7C��-�d:|'+�"�ɟ����\=��x:�B��P3FFo��k��Ǩ��X�<����`?k⯺�hUYt�{����R�P�o�CDn5���L�0{&N�!\��ȡ��J���,�$���i3�9��^�f���򐣻��KL��L/�S�6$��3�����V����yP"�(�F�PE|���h�n4�J:Ի��sņ���06㈃F��ms�X��=��[�k������$GB�f�ªun
t)�
;Q`A-h��/i�6�fO���	���{��8~��F����H;���W�]��p�?���6^@	{#�U�,��I.l�T^e�>-i��� �#�B �IZjl.�D����a����81.����$�A����!��LVy��v����P��y1K���^<��7{��aLa>q5�dz��Q>c���<	R�f� 3�e@�����y0�}��^Z��Gv������=k}�7(V�T����=PV��ب�Q��\⠼I����(m�N�O��f.��V�������+�C�9�@xDB����^�����?�D�G���@�@�ü�P�5dp�P��r�����wgj�R�����r���%O�X��'j�A��K]�,{0�Q(Pv]�2Q���e�5O����eE�07�UW� h�q�I][��)��G�s�2I�9�j�>�VSxdhx��z3 +Z ��u'��@QB�RO�H�C��)�&��������є{�xU��Ua�*��LC�?8�X���5�)b�I�R�ݭ�%*J�/wL�ҍx��|���m�r_��u$S�I��(a�^$6RW��c�GW&:���R$�Ï1���oC���qR9k��D����B�o,�PVO(�G�sI�r<��rp��Y��d	k
��t3&E'�������瑃W���u�է'��c�X�u�nW�7�&i�����Q�� <,N��&1����8�Wu$3�1�cA݂�� 3q��4i�6pp�X{��c�  ��4>��������A���^"�>�I�HG����b薦Sr�oOh���C}�qi�^xK��O�|j�g�dqpgb;�ZD�dp��ePçmEVuU33��Z"L=���B@}��JA�n��&�{�7��' ��y�w覹7������fv�f�1�J�;���/�G�1��~
E
N�A��H�5���d���da��������������a-N�������2IV��	���O��B�!�D4��d��ӖҳΝ}�3�T�ø��|?$��r$n��`�x����Z-^�5լ���ٯ�����P%����&��������l?�q\��
�,hT����B\nwUGΤ��z�K{K�E�X�K�TB� ��	�⤥>�p��e�%��$�;[���h>����?$Z���޲�|鏣2�ϗ�T�mP֍�i.�	����l��ƕH�w�;gn���*K�t��-����B��S���mw�N��<)�;j�{��Z��z[b����"���G	���8�E���0?ɜ��AsW�¿$(�H�P]C�\�D����RBɟ�z��^�{<�#�M�@���Fp�~����^,Z�r5�HݸuS1J����5:4I�(�3���ٷE�����H��7�:M&��z2f�=�)y������A,n�fnPA\7���4�ި�Q~��	D�U���᪗�򃋱�~���#l�^���mj���� �5$芝���im�]�r�����P�lee��	�1l��������q���>�`M�d�Sb`�b(��p\����G��mE��0��k���������`�Xc�L��R���haE���8_���S�=��5NߌIi�F��( ]�-��]0v����2EYԬ�- fCvH�w�B{蚜T�6�pA��T�`m���������\�đ9�R8nϯ旱ő�|UgESi���½2B�l�7b�?P��S��%�j��>@l�c�/�h��'�sS	H�2�_,�p،�٨
�����rAW�>g"��M�a�� p��Y�dx`�ˬ4�uо9�f6��R=��?W�I~;p�C$d`(��X�p);�>��!rt���[;�Wt�ժ���
��<����JO�*�c��8'S��"�=�h����0T*]�k�5`b2�5PI�9Y�B ���.�c��� ,�0d��՟uo�8�u{Ru�?�嘚b�H�,l��Q�q��0*��p�u��-����)nPK#$%g�`�]�jl��4~ ��?�%E,)�Ā¥ �yiE2�A��+xA{z�f����Q�ӵ�=�j;�)��F��q�~L�P�� o+�C̆`_'Sꖕ���yG�[n�Wz�w�De�����a/0���N2�o0L��c�fI�
��~�{]�|�01z����Z���� Ά���.�v� ��C�N>!}L��+~x����:7J���[�$��ր��U#�S7��vp�#�P�@��_�����Ҩ|`u���]�'�Q��l\����� T(�O��C��+De��r'�vʅ�}p�4 ,_եN�7�z�1�P?[JO��o��߀/�޺̬�m���|@�M�W���7(e�0�K�{�)ۭ��F�a��M�����@�,*��eX�AP3�&��HR��
O�)�Y)�\�r�͚��F�n[�y]We��t��)�vk����S�$I4�@�c
9яa�-��������i�m�b>*�կE���y����g��y��3�Qy�R� 6����Q)3h0F��8N���;�ЈK�7dư��B���45���b:0*��J��=3��0~�:���\�b,(�KX�?�2��ւ���=�V������6$���\o�U��@r��� ���k�c8*�Tw�*[� b����M�ݤRݎ�C˽�Ӈ�A*~�G�Wp���z ���7R�K롽�b�'��t'�b~H�V��K �-�|�P�X)HI�G���ː>r�K�x�0K�]r!'���f��[���Z�E�%쀫7e�����-�i����`�1[���k�؁�qgÎ�?�C|��? �۱��j�{�}1�W�w�����mǿ�]�71�c�3�e��|[v���	xy��v8�]lс��/�k�q�#w~�����֏�X'�9����޺�y/���~! �M�Җɩ[D��҄�f�mMWZ���d4�0�	l
{	�V,Ѓ��P�4j�K�YDo���W*J�Y�Z5�L���s	�0z>��&��Sh9�~K���Z���~�TgM֠�(Hx7��S��)��� +EϥDd`G��V���<�z���~�A����Ё����b;!�A�2Nٱ�;��L�r����R�������qV�,&:Q����kdr�����]�N��ܳ��B�/���B��Ƃ ��{�w|&�ܷ���i����SA������u���ٓ�r&c�%7���bVq�A�ſ����a���?UgF����.'�ZDP�t�ȡ���E8�Ӷ�I�_o8��8V��u�
���!�Z>j�����A@��$���� �K0�W�lo[i�Y��H醶�&2_$#pnH���1�N*V��N^��{i��t�i�ȱE?�>0�]_\�A��:,�V�w�sSN3�d�yxj���Z�I�m��C3I�\�ҽ^�E�ޘ�[ҡ�>��?�>�O��{?2�X]�y9���n������<�����r���~��˜k~��Q�0����[W!a�V�tp�)�oS?�p"}w���\E}�)�{��@1�m������!�~���5F���F�ʷT֧���]ʵ�_�H,�*㰳���N�{L���zK;=K�^L�[ݛ0;�e���Tqo�d����j�w�P��/��%E!B�P�>�R���L���Q��>��7�-�ϴ��T&�w��޷��8�D<�Ւ�0��s�14d��9]�J�+��s� �|1|
P��)A}��U�Ͻ�_��؜O�0�e�#}��D��ueڭS���u�i!�i�)�Y�ˑ"�­d2�Fps�5�?�$������%-t��$M-d}1Dg]$��a��Ν�%X[��v/����y�;��xV:���M5O.X����sÅmn8�.M����/�joHL�S���v��D�J��R�t+5%T�^2�'�q��U��e���i�ĕ���~@c93dr�bE���s�s��q�2#�ZӮ�Jf�������1��M��U�WR�֣�/��6鄱R�`�-�ߧ�g�w����
���M�2V�5��Iړ�w�i�A4���"��=�V[�W���=R�S�B�1J��$7�y�N�I������X��9MT��F:oC.��Tt+-�]>�0�nwE����~���+9
d��<܆�/M8�ա;�A>׷hp�Tjc}�������h�uT2�V���N�̛�{�%Ĕ z�X[[^v�����ʧ��FG�}��5�[�b�o�ޔ"�n�joT�<�h���/���ov���01��:� 3�@F�2�7���M���9�Hr���-G��R�����w#���M�,����m���ݧC@u�{@��Z8}��(`j���<����v��\+�h�E��<:!75�J��n0�ڊ��y]M�7-���LG8�tz��3�S�e�&���ŧ�/f��S�Ԃ�N���i'�l�#ܼ�D�A�8K1�ek����q�h�ۋXa>��Tɐ�Al�z{8eF��/}q?�Us�����4�	��5�ʅ��RK���k c詋�	�v�/������r�)SwOl_���`�.��.(E&���&OLhz��3ܖ`k�M�-��~CQD������]� �9Tg��mFTN|�$�W���b���Ǖ�[����L%�D��'w࿿��������κ�YkwQWO��7I��?e�/��`�{TS�~iݪI�馄4�1Y5J�W�y$�|D+S��;�XD!E�����ɜ�_TXM���N\t�7<�d�BC����]_�8��E��*�~�4���������%��N��-1A:Ɗ����?{�lSW	�7~@�C�V)��2Ye�֗V2*��#�K������xnv\S�����Fs�b�R�k}�����k�ֶ��#7���/%۝�)ZiM�l&ͤD�j$v�#����ht�u���n3��w�=D�a�(��i1�bR|*�*�29e�7s@~y2�͵��`}���=a��A����4.a�Y��*$׽=�Ox,R]#��"����z����WwI[ ��&�qf�y�H%+�Vvn匜�#]��/<� ��H4�"eH��y�4 �H���ug���^{��|�E`��6�n�(s�j��^�rw� ���'.^+�%s�46���L[x(����s9S2/���Xfp�X��`�ؽ�q��N=N��]�0����X?U'J�<߯(zI�M"�T�������@{�nx�����]����[��5�|�X�>�>Y�R�4��P�w�J�;[�@MA	W��&	����`�$VJ���z�0��&8���\kI���W�x�j,�@�(�Ln�/!���ԯ�`�!:Q� t���Fx���0Ӫ�>���e�NY����F�K��%0�-�p{Z��_Y;rT�G0{BQ0w3&�Z�N���+
�]c��u P��Y|m�sA�+ɢ�G���Hs<�4�`��Cr����\v�qνФv�-TRo�& 0�ʒ����%�#Cܲ�
!X �ZG	�5-�u��C��90ܐ(dF�XkL�J]􍜢oo�x	�J�[r8� ����ݱagd S�+�3w�s�y-�pn���r��v-��\�l�7�W~�#��wUker��N�.�x1~=�f\�� B�5���3�[���oK�X(�~���+3x�z6��o���G�̳���\�� �9���<\�9�+r�Kb�lT>��v�� R�-f+�G�`�TdE%4fε��~�.��5��}P�e�,�K"���=Cs1�H#�A��ޝ�����[L/HE������Q]Z&D���ϲaU7^F���S��1�]�{��!�h�'v�B�uȌo��W�6(�F4�|xm����b��kI[4j��}H��ʈ��yiH)�3�����?N{u�Y4X���2�--�77CJPM-��^����=�/�X5!-�`'�V�m§ ��7e(h�����&7��#�U|�F	�P�0�ݿ:��:�R'u -�YD�rU��ޝ,R7�
��kD��lr�E��]]E�Ga4�3u�k3s�� ח	�zH=pH�����c|�d���dc���K{�9�.N�N��
�]�=F�������i�8�U�߽�Զ/{j^ҍ_.�.S!T��L��K��Y��bj��~Y
��I~��'�p4��d�(.��Xi#�HOh�n��s�Ɲ;"�?�dn]�(5̄��ep\�x:	�gMo�q��p�zG������Y���RՓ�?�Ba~ |��Έ�r��G�u�>�FK��FI��Ȍ�*)��� ��c4�+���c,�ihR����HSoT��1H��Q�}9x?�l�ic��Ǩ�k�X��^rQ�׷�8�BF�[x+���p�*f �u�<+:}{&%�T���\`<odp�;_8�f�2s"�EQ_�f)��i��V��,�u;1�a���W̛�j]R��?���<�i�Vgɻ�=��un$!�c!��v�аub3˩�>�q߅�&��Y�TEB�P�Ro����R�B�}���=F�a�]X��$Y���,�RR�K����X3��� -Y�%y���/X@�|�b"\ȃGݠ��z��qf�	C�u���S��!�U�~�td�#��\	���5۠ѹk����	���n������ؖ�ۑ=�2���©[�M���%��}�xO +-,����_�aVR�Dݪ��卜9=��܉�XE�4���<�X��bP_�4��!�� r����P�U&%�� M�ι�]H�'iZ�M>�e֪�((����]P�x�D�sHS�
R��Ҙc%w?�%h,ka(|��?i��U�����ӼoU�)�f�2����� D����+���g��D��M�gȔX�@$�Vӑ�k��Wc��s��J�5W����`��_�����D���ѓy�0B�V�ѷzNcAö��
�����M����p�2���剆���gߢT���hcp��Wv@U��9EY�S��đ��<��s�Sp<ܨ�{�7o~��6�ǭ`�����f�O覐3��HaH�a�yn?<B�z�Ӵ��#�,l�D��Dw4yq�@�b��f{F�������k�3j�R_@1��4�����%��[�� nM��sFiWO�.B�S)�354���I�x�*S[�@���e9�KXd�&�R�h��+������by�s-#f����y^P|���}-X�y�B�>�x�z	UUC��	Ss�u�H4�����R�����ʨ�nv���#�@��tq�鸗���I��	hO��0y�{�46���I�_'�4��L�جd�&�|+�Ȓ1�N��+Q^���v@���F��
��ÙŁ�n��n��ٓ���,�|Xa{Z�28��m��H�D8�⯝zU-��`YD�&�	(B�]\��z�W��^̱clШ�X�6��bk��.�#�3*1���U�s�ԊJŤ��h�DX��<�����Q&T2b!�\K5k�x��)�ӯ�
[�a�dp�a�."��vOVa��~�*`�^ɇu�FFV`sN��@�Sߣ�* ǽ֥�O��FФ��=����c���uU�ᄓ�#�d�2H$�� 1���N�?�B��L����F��C��a]N`���I:��v��Ĝ�4�EL��E�`o��=,�ݼ�M���H�q:m��e瀩�PU��1k���:�!N]D?�ݔ���n�Dq�Կ35��8\����l�0N�Atg4��볹��u��ǙqC���^�$��44\y���v��rqQ��gFv��Џ�>%�D�Jz3`7m�-�_��ң�N�GE�B�f��]���f��͘�-P�^�an�y}՗ac�McG�_C��E�;�|}凒��Nh��Ҫ���J��:@�������%�ȓ�w�!q�X�2$��w��d��ozb���9�(Y�}"ø�dx�����k č\#_��y�4�dUIь]L�O%R�ᑁA��Ȯ�~�����.H
���g9��L��J���>�N(�<A��Ѽp�S�uH#��O�?������H����,X�Y���f}6进F]�AhLA1T�ME����4ꈏ����L��w����4�I� ��Q8,��0W�YG�7������sӎ��K��v��co�M��0�����3��G^��9�/=4��N���1��3aUD�	�b�D~r��
J:P�nզ��o�s[�r���-��CH���� =��R��ߥ%���(�Y�e�x�� �2�S��q��&��5�f�Y0�n��҆����妖,�Ֆ:qCR`n�Vɐ�^W�8Q�}Á\�����޷�΁�^���������u�EsxGFRs�ҫ��C�(��$j� �/ܣ^3H�4��$�#$l')����0�A��#��	ԇTo�N���������ȧh ��T �s1���e(����m`�� �_z!FS��V�<1��>C�\�8�'�R������~�C�-� �n�荲���Qֈ��[���� ����uٴ<�d�-[���~p'"��
1m�݇X����W$�:p�Z�*B0��T�s1L<�k?�p��6�x�:\=G���&zk�����e N!M!�!������`p���+t)��f����.�)b	�	<6��T0?�Qф��\5i"9 ���]Y�hu�����JrH��2����=�ڽ�����O���=L:�}1#^?�#��k�:5�*�
<����W�'�N�F���%�{'��������"��oB๨�H��B˺{��A,��-DN_��.�[�^�F��6� �-g�L��M��b�Dt��h��i��{4�濦7@1�t1���s��'���E\�7��'�)W� �Պ2�R.��s�M!�#������T�S�SyY�ꢅ;�\�Rlj�IP>S,��+e�a���c�m�te��'�B�ƈ�g�C�E�`��^7�J�?�B��oF���ٿ�6�bR�w����ڠB?D��M!� �ݙ�-��(��?�(�!���r�h�� �מ�x�.�X�RQ�P�[{-;�pj�K�0+OY�����ǻ��N��wN��ӛv�w�J���I�B��=�*�F=���v@������F�1��}�w�2����:n��ItED�v�x�G�ctwz��9+^h�a�.B���Cϼ8���X�2W�4��NK9 ��R�����x�N��vvA}����
�K�1��f�C���+���WQ�A(�#'V��/��X�@�)\��:,��`��OEj?n����qLOSS�&�S�l?��5��>��0D��Vq�Ⱥ��oV�up?�`�3׹]���K�^L��� � J�"Z��R=��W�9#�s��Fx�V6uE�h"]�{ h~F�_á��TŤ��k��/�Y��=hb���o�w26�t$:�g���SD��ض��ۖ �!�pu��e���ڃ�GUp�ܤ�O��ٴTυSYE�F����dp�q(9����ރR��Emu7��x��%рG���j��s�<���E!1�/#�p8qy�B%*3�`vF&�pv��ا����U|�}Yxqa�3�3eԊ��r�d;������+��}������R!|HH�
G^��i�h@}�t�m���47����L�l�� ɕސ*u�nc
�����p1��lB|]��C�]�l��rn�.���ٜ]J���A�Z.�bP�8.�X&� G1·1G�Q�9��l9�w�y��e�����L�� ]�
�X�Cs/�X�Z�H�_C+HUȀ��QkW����'�,����ɟ����P��Z�MGY
��⯓-�#|��3�D�88�'֏z4�Y��R�6���Xc�g��I�D"-��*�<^M%��V�Ɓ�4Cě�� [�Ó����%E���P�a��d�����`?<��Pn��T����W�+2%%��R%~ 厨�������1Y+n�S%�a��pK��O�����F�b�	����jJa�A�ZG~���L?L��|���˧�@�h~I���Aq���i�T�:zUŭ+���i}�W�M�=�P���	̤���iC��)1�����Yٝ5g����2����1<V����昉G�����2��p/-p�.���(�r"���:��0R��3v�Ko�t)��'�V3]W���gX�7Ph��1�~�8�N Ŋ�� �ۓv�W��	��U�����S"�xD�兯ʮ�ڠKu��
����{�j�x�O��Co��Q����M_�1�-6̶��֤�� �x�f�b(#,`�s�a�Fq�zn0~�X������P���P���H`��aq��h�:k��	6��*
�(%�1�P���B�4v���R�:��3�U�j>��EH�����& )��\"����I� pLBMT���]�������{�ë<�@���HRq�]�4����^���7��`l1��"��P��ѐ>8�@����Og�K�^. f��	���I�/SphZ�q�}���GÎ@�4(�t�* æK	H�p�ی��jrG��:ʷ�|��"hoD�<��)B�Ӎ���xdǤ�!8&k��UM�Ly��q���KĊ����8�]Wuv^����JQ�z��@���	�L�h���}�h��o?u}��{�6��T~��-ozi���/��Q�(�N�W��u��޸x�o��/��h��u��N�_S��k^�6��;~��R�O�+�*��c6�áے�9�d��'UR���Oz���Y_���Չ0S�y_��s]ßc�s���Hw��t��~�2`�JY��ß�͢�bцݫ`��@�����]�g����l�\�چ�)�M%����Qd+�Y�RVʂm��L�Xh��T��	���1Sd���n�k������GT�}[� ��^��ꠋz�s䅟_غ�.z��o����SP��V�;�j�!����X�S��Y�k��z$��N��`a�mY��/~>�u5y��w$8e����K���:�T�O�-,�N����wB�F����~2�鍸�@5�9�z�MVu*.z�¦��,:��
�:z���\��Dt�ʶ�ia�B�)��S3�Ҩ�a@丹la����n0����Z�󌴐*�����%����ǋ�z��T$�ͪ(L�2�����w��s��2��7�w�G�nB��q�����>r0�7[4�2X�GUW�^H!K�`�_��������<���fk[Ϲ#��/��yL!Z��H�u�
�$^
��LTg��H0��n[p���:�:xR���;��~�FUF�]���3*H4���hx^���~��i-5���K��f�v�p`i�B	�&���Պ�h�OM���ůص�rPo���#hj�n!���ܡ��m'�V��?(O
#�R�n�8�b�� � u��� �73Ky�o�Z���PyL2p!d;��� �L�w��ᾊ4њb�ډ��Z�H��ZҺ�,��
��$�$x'E����p�S�����~~����?c�Xq��Xf:ڂ�� o^Ն��~
��L�{��ܖ���<�+��p�E�d��đ���� �P:S�;�Z@Dq[�Hy�.���87Cc̈�v$*�]s[�����H��d؟�QEAjW��q��S)S\�_�k)�@��9T��%�9�3W�r9ڋ�p����:��6��IrG��c����*��Q�PC�`�*��Xj�6y�=�ȉ��^�cp�����S�-�ʴ�&�L
���4I�;|?`"�k:��
ӱ�k��Fvj�	'h�ߜ�oJ�I.�:���B2YR�ݶ�韐d�1��%���d^���문s`�KJ>�;^�x���?�'�@��첝9\2�B	�����s�k�^�g��`&N�/����Y�kBQ�\ �	=b��3�T[���2b�#���~���0�V�ï;��w#�v`c}oa��k
�R\zK"g��L2vK�Ա��&9Pw�X3Q4T�S��_u6����L�����f�-������,C���6BxyǲNm��gF	�f��L���&E�o�����c��ܾ��֟�jUT��R�K�)��ۈ��<C���d��Xp�o��ߐ"�2Z��.�F=�<������	7k8�&2l���~)�L���<�8�z�����T��#��Me�P���
�C�L\g�%0��!dr�gݜ@B�w[�^L�V�P��g~�~�-*a!�Jz������L��p.A!��S��ט��ԕ���a�]$���Ϣ�2Kc����yt�{�E;���F��)�~���z���Ҷ�G��-eCH�4�kv)�v�Ȓ+%L↏Z�o��G�[��G���t�Z��\+��5�ؖ��oȾ9�/it�~��F��KuT�`�%�i�+��#c���W��ʢ�sO�h� �d�2�1�!DB(�.7#�W+�7DqU�oġlrHFa}"�J�8�﨨E�6�`� G�/M0�E��2�����a^s\�{e`S1܃���!!��P���[�M������.$^`X���K�6�"�I=���u-]�8��l��o��c������3����>����4�_	��K;vPX٤�﨏q���|�K����M>5��r��.<�_�|�%n�mz�[�b�����{�8.)�_Ysfz�<10� �����p�V\mHݻL�½g�Y�&����>]�7(���(2�ih!���$:I&��mPc8��/��I��v������K�1K`�I�z.+��n���÷ޛ�=�G T���9�\P�Dq�,k�>��!��B5�D���T��QmŊ̈�o�B�<�o�����-�s�U(g�I<���Vⷎ�;����эc�rF`���ix�|&|�1����R|���LG_謙{���	���+B��@��b#=��㇪ͅ��Lk��)�x��l���I
�.+��G�1�\�YU���pfڡ��I�&(�K��φ�R��-�Lzeһ���p$֧d�%0����[��H�>=����`fI� �� ��7�B�
�L�_�&_+q�I��\�R�L0���v��׍�:|ڌ����<�B�9�]�?U��F��EF�����Q\���u9�*�u���m�
�TWʭTb��[2i]׫�&�?0�������WBŃ7D\�$������s��!P�Yb�}ԊE��⤌
�)�-��B���Y�f���E���� [5�1|<7�%�r�s��,�����ք��������PL�}��������O��'�C�K�P=��r��~̆��X�X��n����T{�#�_�B�A�����;0���=Hr�`})�7c~�DM}n��iRE:�K�ި|��������RQ@9��j����1�/�g�uu�ζMR!j��<��+1$i�{O:���F#_��TM�a2+���C(���a�n���zTp�}���+�sJp�SM�R	���q��I\�jP��$  }9��Ҧ�c@��Y��q���a{��Ұ˙=Ykc�?D�	�%{<���"�f( S=r,4t�7��fX� ��^AG��T�}\��R�*�_�N�����@nՄ��N�҉?>�/�q=�%�ހ���q��m ��L��}�ɥ��Y6ds��*.J#[f
Ԗ8�X$�ߵ;p
��nd���yf�y��Kf#S�"*}#��"YS��M��$ҵ�bS~⼠.�B�R��z�zf��r��-b*,sB����L���ثڂ�C�mФ�$�֝�r�h��f���N9������j��_���:�XS���/�<���S��!�:�����޲�є�e�a�:x��P7�������z5��*�!
���^�4��$�>��a��!kNh��g�ffT�S}5al7sѰ��# ��ڤ�;�aI F��T=<��uP��f�k���l�&ϋ�Ǵ%',y��K�#Ϩ�BQ$S�l��u���L��c��9?��Ѥ�{�V6�|ũ}a>��,�q^Ym��?>Z�뼓S`Z��L�ˎ�����M���^���3.���:��?�+9	lڔ�*��f^�	i��ů[	[ݨԱ|�׹�JG�,��̀M1j��ʛ]�t(BM� Fj�����E	��}.�0a��5x�(Rf>�����%`6Pe�#�z��pF�O;C�Hw�5kԷV4Zy8$�i08Ӏ����O��G)5N���Hy�	!�<@��4*�H�.�Q%�s��Z�%V��fhEaξF��/ڏ��l�3d�Վ����&�ދ�8���`�EΕ�c��s�,�#�5��6@�#c�!��*�b{>EF4|��֛)�T����}w>���	����?~���;��*�b���ۼ{h����yj2��!��U�����6���#8�Y�C��I�_�[c��W���M
A� �m��p�66B�Fc�M4�X[Vm�XH\����D�L�+��&S�p�����d.#Ӱv)�Ta˷Ǉt�lt��e��8�|�B��a>}B�����cFt��C~ �]�A=�6��Z���[���/C��C��=)�h]2J��P�ᗖ��R��C�?;ĺ�i��A�� Y_��V�/���a��#�̩_0����H�c|�O`�Q\	��L��#M����qB��q)[�ߒ�U5z�}N�WM����������k�m�gT1�z��vJ�G�ޏsh��R2���M��8ǚgX��2L��/6��[k��AПb�w�V���֪$N�w�q읽�ɧ��{��E?W[�s���2�6���ׅ�S�m�e��k\���A���Ĉ_{����������L=Y�_ʚv������0�K$A`ny�T��](r	O@�/�EG�^���4���`;�Wn�M��N��	|Ze��)�"��Y�:�5IT,@�y/�8Ju��[B���/�ϰľ�*�_|y%D�o��Eyf2���3>[�Y,�k����?���E@�G���=��(r� �!�1�K���c�v�d�ŕ��� ��X��SEV*�m*4��~ߦ�-����<+�������t�|%��Y��Ć'/qӼ[ٗ��@:g�uXb�cr�^ m^,�N@e�-�0����N���O�i2��D
LV_���{���- ���n�m��M��4�ϕ�(��Bƴ�I�l ����s�M��r�o\S��ψ�/Ap�3����������&�"@[��ȕ��۽�!��n��T���+r�y�E ~�»8�mi�JJ�V.K��*ɵn8��o�ӧܸd9�#��k�C+��j6F�:�����>N ��J(q�	ǘ��Ҏ���~#`�Z���+�Z��8V��d^5�D���2�#�SW��|0�\�c�pe9�������v��wܑ�����\�&q"a�6sM�Z��w+�F��Ϯ��2����b�B)��HgJ%��#���ۀ^�B}�7��e2 ����(�{�e����5���2l����-�a�4�1�s��=��#��+��,�����lb�d)W���z��b8*L�[������B�ԟ�?:;+߻-n6�N�J���(�����־��ɦ���t���^1��Z�����6�׼E��P�����j#������f� �ڷ�������3{�.M��Kz&��[��;_~�Z�Ȕ�%<��hpmQ�]f��(��(�30(�vU}}/H�W�������%�c7��m[Ƥ���9>�b� ɨ��G�IIvw���\Er�CEd�Rm`��9�W`�<�k��h��B�O�������e��pZ[.0��ګ��p�/Vk.mb�<f���ޖ�T!�o\�;�Ba�4��"`��W��К���2�,p�K�����MZ/��`��I-V�^�l1!�0qk$h$=@#%�� ��\0UpC��N��a�W^l��"(���j�}�@2g���~I�֗+��v�Ax�Źl�L�)�yv-243��42j6ΰ�]@�J��
�K���:����,������vc���#��F\�||��@�Q���O�<Y�G�o���ק3�r��jnd'˿���ڿ�5��?����S
��w� ]!%��.j�#���1P���?�F�Von�QƠ�ƽ<��A�X�פr�&�K��/��9�Ӂs���؜v.�D�H80'���e��~�¦��uƸ[�w@Q�����[*����ԍ��o�R=sf�$"�ʌ%-i�~<}�k��mk���4#��>�s���	I�����|�M��;�w�>���f̵�����MS�#����r��m���0��S��U��M��i;e�	�G��P�E�Iq��Q^+�&#'�SV�	A&7u��_S���K�����b�pC{U�Ј������g|����2{��B`��G��7�k�3���[H�<A](�]��fi80���2@z� �~S!��
V���$n��Y��NP�t`�"�}0)�n��Y;�Ca!]��H�B��,l��sW�Lr}�Ɲ��{�y�3�NcFxM�;�(���Y]p�zwh|�".c�?�u+KtY-�?u�߬�-���)�Pn�ǹr�[�mq*>��!T~a��g����i^y�QCۅ��ٝ��N:?/w2��O��U+/vw~�}�k ��O�_n����q����<��UM-�\:;���_��W�>��������=Qv�1�ؙ�h4 �?٘:XLZb�1�k[q(h�:�t��ݮN+���@�#e%��8�?��HH��z*�d.���U �i�=���������j�V^މ�[W���?bT۝٪m�/p�ɉ�ץ��-T��&�WŌ�����I w<�&)M�c�K�����j�l./�C�A�Q�����Zhp �����PL�������Gvz��� N� 9흙-�G�܍IQf�8�W���C�|B4qe��H��E��
�J"��T��]��BG:�%3�����b���a���v��a<&��B"�)"�^(CM��70�
;�}Хf��[ś��釒�~ܖ�c���O�`�s�ȤAq�\�\BWN\��w*^�Q!��|���1:�%����M��B�ݑ���=r){N6����BwӃ}��!��C\\������&��r�
��\1՚�Y-�?s`s4{ �3���J[2	@��w��|`X�������UZ�����)9A+dvUM���Fi��lԖ�A�l�2<�	3�@H,��J ��,}l��M�U���v%�7<����Bs�ĹX7w	F��k"�AO!���X�`]�����o
��*);B5r�D�ӔqdX�õ��f������\���ȑ����9z�Z�V;fs�`��ȳ�ģn�Y��V���,�*��Z��}�~���@[S�h�*�AE���Ƽ[��Ld4�Fl0.���/9|o�T] !� `/��|y�	j�z{��{.�'�����~�������(�&�ܱ�Z��-����/Lv&��\4��������� {�s�I��"�@�<�A��v.��=\i�����M�%��{��=�[0GI�c�$�~@�5Z��1i�-��`~�tV�U�_���b�P�I�-!�h�B1N֋3�(2��cc2��cB�%� M��R0���c��om�]��� �S|���Ş��¡�+_�� �<�^C�ڗ�`T��;�uC��T;q���L񝍗w�<Y޹`�y�Aƽ��z[�����7+s����I�"5�=]N����q�?��ɜ��u��x��}`Z�[��f.��&�SǸo�`
�Ǥ��9�I�P�>�ah���i�D��Z�L٘��u����~; �MAǑ���,DY��|�2��[���E�7,J. �|�[�}�K��Y̎/@*<I��b�����u+k'�Wc��W+vX�';h5 Ȑ	���ұ�Y)Q9K�Iz���k(���Ȋ���Iw���g0A�
*��OTx��!A�-P�[���N�e =
 ���<O�+t�	
�A팼ڗ��bБ�U�c���Q�=2�$)[��k}e>̦g4�aF�%��jo�=�'h(��&,���]�K�d(؁��A���0	]�2�߇>��S3f$4Pf�.};�����ġEo��M�O~���¯��J��#&ܕ*��~�-�zONF����Az	����2�E���ԩ�-��&#�J�5���q[-��NAެ���iZ�=s�����ch���3��;�u��P�C7�W,��,��(��f�;�J̯�I�<��9���'��(�KjS%�;�9���=aQ�8��!�u��� ��]l���S��E���F��-�c����}gtUS��a�qH\�vZ�BZt�fE,4~�MۂIc��W-_^�U�<��M1{�CB������n�v��_�>9Af[������W���@$ʓ!���2{'P�<<؇����j�7��$N�VM��o%HH�1����	��g}"�<��.���\lS��1I����LE�S���AA���ij^���%��'�e�I��=�LRΥN��M�[����G��.\ck=F�G��������rM�'v�J�t٫u����[�W�q,�� ��|�l҃����U��>S�AN���� k�(-�������bB4�x�I��c�)����[ů��o�;�Ӎ��HI�2zͅ��:3��5xB7�w����.�b��s3K����}[�����K��MP2��٨�Q?�z׿}�Gw��={������3Zd#*_�5�y6�� :`tkYnN���;U߬I��l���p~E�(hz�H�1����=E���:@╭�"�X��M�"����=߱��^f�s�ޔ�U�*�ζ�(��^V9�0v+�F�_�'� Lo
c�Rw�B?]�9�)�����TB�������q�l�,d6�7��<7w� ��_?�+�#4�f�Ʈ��'G�F��֛h�FPPf��%F4�'>�7� S7�2T-�aXu�ѥ�?�cק���-֍�Q`8���1�M��2�G�ûe?Q��Dw�8D����gV�L��)�8��܋��2t󷼩Pz=�d�|�؜��'���6�Φ�����O�.Oo{M�ƁOkR��Mĳ�F��F<�(MaQ����:�:LJ�M!�����6�A��}��.��5W����*`P�W�KM�8�Ӛ;����b)�D'�S���
���h����_-E�!�
�"�"+Zj�Ae��?6oA.g:.4-������R ����`�Q��)��X�����ϥ�2����"i��0��Hd+z�2R��;�$��T����10��0��N�����9��{fT���Ñ��(=y*����%&'J�oC��%G�gw����ώ)j�n�5�u��&ogY�\ hlFb��k@��\��+~#���jv�,�l�Iz��<��?�}��nϚ�X^�7��h�O߳�N?;TX<^>z�Q�C�jN6R�i��Z�p�=���E�ɐ8T��&Xy*{��Q:�?���(H㡙���g�*�<��#��0�D����t��/j�%C������C��HmX�V� P�Y��d�% L���}�Zr���cM�i���Ȋ�}��\��l�r��P�7��m�"��zs˥
jz��}�ER��M���I�o�!͉vz-w<�!;;��I��Y��l����4>Iێ�V�v�ɜv[
%.���n���<�FGF"�k`�%m3 H.l*F�5�䧱 �p���|S�w]~N_c[�Dl�`��w��C�Rl~k������0bgiy���C�]�ǟ�k��L�׭�S[��Y�c�s��y��E^�w���cP�S�z/�G|��8�Ca�f�_#Q��T�����$�2�`��oz�O�Bɵ�͢�����Wlf~R�^��u��-R�܍���Y]&/�l��̱/�#��I�TF&#��֍�Ap�9���� �_�ĩ{�呫������I��-��\ժkٛ��c?���~*B=oH�]�ʃ5? ���������8̑�5!��2��b���&�fY�k7��χj'��f}�}�JG%qAT��JurӰ��6%j���F@�r�.�.v�eO��
Pڅ�7�k-�h{�{mͳ4v.���?���2����`�eat�K%-���p¹�z��8� ����gcܹ��z'4^j�9�2B|��I�VD!��|2��&0�7."��<�	%r�2j��N�eC�M�5zMg����tFK��5,�6�'��dv?��+�q(��b���4��`ih�qq��xW�fF��/��8��R$�	�t�_]��+x��A����i�e��]y~�ZW�x���IR�0�,>�h�����#�v�<�56-��e��"@�F+�]��q�=z��X�M-_��5��*�9�_M����b�dN��bb#����mEr����b�b?4L"�@Y" '��'՛��_�1�� Z_�3�ţ���0[��B֎�^�/�ڽ��?�Rw��
9-yr[��:	����I��ߐ���c$�BN܋���<A��C��!=���4��C�^��We�E�A��U�O��3��̻�����}�YJu@֥
���t(e��2���8H2���)l�����m~Js��9�N����ϻ\��U�h��&йť�$0S���a�Ohi����t�JJC&�����7������q�s��N4N��!|GLJ�8[T���KE��c��#Y/��ؤ;��*Ux�l~���*W)�'("��AY���R�49���~B�@�ى)�H�s��ϢY!�Yo`�$������3x�i)sW\�x�u���`�]�Ce�!�\���Q���e�D1�f����}��,G�p�^�ɡsǧ�}1�t���/��]xG8R������(�j��]�Z�^o}X����^��!y��M��'��$�aڐ���S{/J?��E��k��y�o�jŪ&�.T���2@&L�I���F��p�twZ�O��9,t�ap�M�Sk�Z��yW�����cL����)�*XX3��k̗�*��[EƘ=�<Ot��m����A��}C���t��u�T�f���y� �i'��I3����HV�H�nS(x��|�?���.z矈�<2�_�T��p� �O�zq�1G���:+�1��c�6W���&(�����Js	�Y}�v:^� &����\���c�m$�L��A�h�W*�1|袏��7��%CT:}D�"���|<S-U>��a�;V!Y����G����caw)�(�L�C��;��B]A���W���?��Ɏ��B��K��4;r:e#�-��%'~	�6.X"�n�rma��I�g��E{��r2J�=�LQ�*'-�I�Pֹd����~er�Ᏽ�s��m��uF}{m�Ʌ��zcO8��H�p�,M�P��[�Z��sܼ�C���t�u�V*��RG%�� I,<bx��u2E�wɎ=Fu�ā�R&.�D�8s�s�ĊX�_���.�a����V��9LEʧ/�~���5��B�_�R
��ޔƬ@a�TIXd
;��-5�h�H`�7~�BP��c��~BY-0k�d�՝nr*V�..�Ț��X��P� ��Qi*�f&�8�(�W]�5��>fw��ݓ�F����` �a}
0M���u�X��O<����g��G�6P��xI+�8.�7�<��N����5��`Q���SSl�q
(��N��;��'c{LQ�>��`�+t,L�~R���j?�g�%���U��S �2������؆��=��ut^�_y�R��J,,GRY��������	})�B�A���BSlɉn\C��K=��0�x��.���Z�������6�,��A�<q�&k[���a�P����Ԧ���Z���s�M<q��z�V��:�q�aP�]�_}m:��nwV/h㔭�g���C�&�gޟ���ct��z>3�-G��dY1�5���6�k�u�N2�(���_���[�^F�e�C���
�'ʐ�!����[ħl�h�CハW&W�������|g3�^S��w��}ጷ#���_�a�Z�;\!k<߬���F`���ʌ��P}�`0r��1139���:|�T�������36���5�܋1����F���>r��bt:�w����o@T�@��n�~�`kry�U؎a��s��
K�^/\�3� �}<g�Ͽ������UF���z��Ŀk�*���m��]��u>r���6��و$K��vF�G��~��F F�'ؚ:PJ������P�M�֬���L3d�6�S�,0�-����1��帼ťwל�B��OZxV,�NR7��x���v��ج�+.��WA�e"���KcR�+Hp�Z�� ��G���V+�j�d�[@Q	��L$$KƁ��w��hI�X�r\|g���ؿ.�(b��J������hrI˽9�����N�g$���	����z�	�Y�CZ��!_��7а�M��B��ۊ(&��Mk�G,C�t��qY,�~ ����SLᱦWS0?���yےc�.絔i#*"��`�7��&����'Җf��JrY ���Ƙ��(��V��Ա�,�b�?����@��$�����T�_@�oʜ̆1�g��ș����wd.$c��K��7󤘥��'�X���JX
�u0Y��]�D��M�g鉤G�	������MgC��M�c���PS��|lQD	�ȳ�����H{�?��7}�`�6���`��B.�edFt�_9v�JC���ؕ���?(���{a���\#�Yo�y����q�W9�ՠ��j�0ڣԒ�#�} ~�w[~{c����R�NK$(���l``�y����g�o4�@aYc݁�ԄN긅=c�m�<o ?S/���B�cf�Hw��e��.C���}��z-J�<��2�ģ֡���V8{�!��&no���@��,Wv���Y�H���j�5с��6x%!��������8���4�YE�>EP5}�����?��3�VJ` y�Ъ=�3�H�_��3��+�Tp�i ��ؕ8n���'PA<7�D�����R�	����ʗ�;�<ۙ�$"^�$Ie#@Rh;�嫑�b�F��q��1�s�&�^�OH\���yP(!�dr�h���G�ΊjZ�h���?������g�X��X�Oȇ��T�й�\�=�YV��5��AH��]h�q�ܩ"Ӕ9-䱮ɋ�)��?��|I�t$F��:���^XǸ"�<�.t���%BB*��#u�.$$	�
?���nh�@�����b!7����@鷗�������g/��H�W��6W�]�D=te�1>Κ��vO����O���*\��I�c�A�2%q_ߟ["���C�Nl\2���h��Y��H��Y-�9��^	J�#���>^\�7��7�oPj)�J���:M��5��#�
�tC��[lk	k!rP���O^J��%�{��Ɇ�[�6I�g؀d�qe��u��ާ�7ކ���lh�[�X��m�h�%V�A���>B������֡��c��q	��$�Mn%���V4��2�c����Mv痱`�u|�$RJ[��0X�	!S��-���|a����-ƿHd	
<��K�q
^����4HQ�t?P���Xw�8:�\ԴȔ��h��d\*�@�4����0ŭ�p���o&���ƺr�Q�Ek՞��'34J;�ȷi��|���[!<������@��Y�FY?ڶ�n<�&�6�y��9)���DGL�%�������H/z�Յ�m�AU�������~���T�f�ʔ�� �,��7�����0aL��-�>}d�=}c����k���L�;c��ѪҨ�;&�H��tC�@�x���\';P����a�����t���l���UFl~g���7���rQ�T���]{����.�N��k�sӽׯ�4w���T{�~03��5���*�����~����rF�F�ê5'�{B�~S�`�7�&wF��
��l�Oѯ���o����)�&G5�LV�_o�v���:�zzU�X<]�Uv/���5���Ǆ�Y\�>x�bVB��q��d�:"��a�a�H!�o�|8�u�z�w��RR���u�������ek�c�YQtZ�)�c�������gvAY�O[S.�a�er3a����z�W��Mr�����4�a�/pg< �W>����}>.cM�5�x�W��r����4���9y)
f5���<�?�����w3em.��ޟn���~ ����f'����qxv���� ���ϰJTGգ��k0Y��@X�r.���^$����P��WT�T���vz�D�9`F(����j�{�b	qE �܀Q��
��Z��-c�����E�ۺ������G�Eϰ�&��3{џ���A����S�%���B��̯jٶ~����8M�(�q�S͟�d��o��.������5�<�)T�����U;�n,���SV?�`�6�9�QJ�`���^G4U*x���-5�ImZ��8u�KK��̳<��\ b4yo�:�I�R�S�>J��RG�M,����D���q�� �k�2��!X��.�*A�л20h<���sW�/�r=)��x��T6�[KQm�}�v��Yx~�$�)�@n�.C{:bi�+,4D�U��Ǿ�Xl��]�>�Uw�o[y��g�k�U^��J.k��(����k<��f�*�j+�R�E^S�E"
K��	]h>>B�ְ��QUA�va=+��d_B0�^��ɕ�1��\)ۄc�٠i5��� 8NC��Kz3)������!rH<�_gn�\r�ߕX�@А��	�ď�{�i~��8��t��%�COE'�W^�Fn�u�t��\�7L�RK5ҷ���_F0��7��<����:v���=`-�.sQ8�$|�"��6�\N�V@����=T�q웃��k�9�o�"��	'G�(g�`{t0���?�����8ё�Zt]r,�>oh@G�:��x�EP�G����Et��R�ĉ�w>Q�;J�^1" �w��?Jq/���<��u��\�kG��h;����p�p2(�:Lj'O�bV2<Ե�B�$�����;9p����/�7繠&�O����C)k����k�L�AG͝�	4�Q�~YIQH��sQ�l<��x�FlAyRLX��Grh��l`^u��I��)�(c�4$��o�8�Hi���֢9.߾9���N"�]�nϳ��Z���i]��hX5��G*�1Dm;�M��R<c����iSa����4��!�3�.�T��W  ڪ_;�H�q]5�cv򉩁j&nF7�Am�gu�@E+zSu!P!�J�TI䨨g��cӾ�d|���B#]��\[���ezq����8��}d	��DS�%;�p��C4�Y?l�:����KB��ªȀ�g�y������7>R90�HR94��ǂ�O�
�ZDB�V�D_�;��9VC��&���:��4�-2������?�\NTeҳ�����4�O��
 a_�q�����L��ǝ�3ʩ���L0�MZ�F���(^;;��u������?M�S���Ш��/'P#�()=������h�	\��i��X)
/��v:����89�Av�R��y�k��A%�@诎`�wa��AC����W��K�}Kp5��i�~sw��
�	ƅ�����H���<4�8���! ]����,�ޔ�m�����%7���Ws9������96Lhi���EG-�E���P�\TA8L�3�3����?��Q��u�����а������H�_ҙ��[D�:e%���)�u�֚N]������N.��+�#��دN����p�O��,ݦ�)x�h�>�O��Jm%m�`��Q�O?H��R�
���G�58�ԕ)�T�GE��E�=u6(#��X���)�V��ZK�H@h�<$��V�z�����"�!@(��v�H#���;����K��8f����\޻��e�G�=�c��NWO�ޭ�qB�]D�E���,���m��ڜ5)��{^�q�fJ]�#�<��x�A �ŤC㷿\l?2�u�"�
a��{�	�CN�fn�8gמkm��V�?�VRb�6,��_w�--LBּ]-UJ��[�����,eA�<��`�I�Ȧ#�SkӅ�m8qXjM?��6���2��Kن�btK<�ϡ%}AXTZA�k��w}��� ��y����
�4dP��7`�����8��&0e��k5	/+j�4˞�V�ʦ4�g����z�!^��a��*��>|j�ZiI�0F�IX�a>v�Հ�4�g�4Y&��xL��2�X��T=�s��h����i���<�L�<8���T��3^:�� �b�%!s0���ӓ�5�H�S���~)
K�y��T 43�Պ `�6�ac[d���6w v�fT�+�F� %ίq�Ȓ'}���J<%�,�O=3y+n8���5gS>�H�����~3�c^�_w"��h/���u��~����oR'��I����J�G�D7��7���f�_��}����i�s�;��J�k�>�yu:"�;2�Y�S	�oo�5�k����|L���Rْ�q�*��P9��ãQ�9�w�z	 �Y�/l�53r�"X�3gc.˒����zo�Sv�]X�P�Uޭ���6�ܒ���o���B������M�wݢ�L���(w�g+��l���K���}-�:�f�}�UC�%��z�Ȏ���[1%#h ���9�U���Q���̕��d�ACdwZ�?� 	�����t"֪{x��=����e�沛�݅�9�Y��k�3�;g]3�x���OI;��m�fEXW&DqO�:&6+ev���SDv��Q_bZOb�<�4S���t��_@�*f��S�q�L�F�!2j 8ʁ)���\�83P3ȵ惝^��ӨW�O	aC�'�����%B��������4�n���	�.��x8$�u?&��3J��� ���V>Ƨg����'�Zp�w��8��}H���v��1?��cF)v56�#�9b5"�ǹ���<� k岃���#+�ӵ��l����]�e��b֪
�a�Á[�6;�(`v�zߡ��F���^�H�G�4�l�ϑ�r�u+uEM�j,�>�f�E����o�إ�T.���ڪ��Soo$r�cs�M�5pR&�'�:��������e+��C�(���'8]/?jS+�8�.�l��j�(���5��z�C����9������t 9��	�k�����m|��>�4TAs���3͌�m\~m�ǢUCqԔ)���)k5��cDg\_Rt��d���׶�2/����ŵ8K����l K/e��I �V���� 2�ψ�H�Ԭ���.�g�u��E�R��Qs�����C����ǖ�䁸L_s�:�`3����.�5��b�ޙ]$r��-1�}��1C������ңǝU�c���'�os�@x��5�S:0g8�;��cݍ�n���,،M�)_1
߷4�dP�y�l!�8醜������"|/�����u�c�����S����q҈��Vԑ�h�����Ϝ�j��ޮF�27s�Õ�L��J�N�0ɻ���R0�d��QLzr�g�O%��
W � ;�QZ���䬈>	��fr!Q������/��Q�R�)����ʠ���}-����������w�ZΙ��{��d��B�����U!�!vR��M짠Ժ�����S�HʆR�����V}C��� eu�xuaJ�Ha�N!!��ʶ�tZ�B��uOd3[Bu��}��	�i9��?��H��q� �0�����`��jE������\`wv[C���3�O�*�4��);:���3��$*G։6n�������?�ɗ��@��;���ެ</;b߄���Y�4�I
���|��?5������-/���S�qR�u=�<K��"N�aO/�������A��/�\�w�c|�X��++�����):Sgi؟m	Nu��:RF�����΅����"�H���� e6�<� ����
���\�x��ᗅb����p��[1L��2�)�y�վuT�޺����O�ߪ�w�5)�s3k��g��ڥ���,;M@>T#��G��F��.	g�	�����'~�y1��1������4�T�y	l���R�G�4�tzT=����y|;���.��Q�M�)�LK�;��M�����O4kj��0��%>&ѵ	� �a�\����!�jz��Э�ߖ�n<H��L�.�Ί~��=�X2�lz6���R�B�(�iӎ��OA~���ͼ�xԉ��u�Wݍm|u�7��4��qF]B�����3K'
�/i��"����J/���)�=����.{����=N���u_.Ч�N~��И�X\�Z�#��9)Ŗ|�]��i$�R���#�0s2�CEd��J�&�Kd<���FL��A�RX���"��5s��^Oѽ�t�T�.l�R�>�]�[�?i����,S�"Z��R��=��3��woS  ��!��`���s[eCh��Y���B�2�F����^uI�TYޫ�E� �R��wv��1���Zۅ��Gk�<�{���mAfr9�����*������|4]��L��s�l�lc��<�6��{z��s<�IzT���ESg�����1��He	�C��/��꼓�Ttd��,w��枠�&��R����G��NroPQ#f�|k�R�m�� A��b�%a�
��`�|����5L�-`�Q��-�t�6�G��4anc���\jf��"��=`��H�b��O�L�g�N����1~�~D���W�Ǖ��15#�ﻜ����u�M�5�5kE罡釙?�������}}/C/���x��I�\s��QFN��;��u��)����J�0x�k�/��_�������ӑI�x�t	���Y��ȆZ������L�<�����1�7��rP9�ՠ	"�����6N�4v[�� �3㝆��G�=/3��>�5��O��k)Nq��V���:Oi��%�jtxƩU�r�ݖ�R���I���5 ��N�3�,�kMͧF[Q�+?@�yr�(�Ds�q#+kSdF����A�L�Oc��u��j�kF�<���4m��ת���ʍ��d�`u܃Q������-�f�҅�v�!z�n�T̃�?�}�CB�Ҫ�դ��F�-�Hr�[!͈�q��lY��^u;Y �72�N\�>ʻ[�5os,l�^-ms���MŗcE0����Wk�Ȼ(YJ�u�Y�����0�,���2���[�aQiC�)�L�ڨ�>�F��(>2:(���I��~���^;=����ZȢ!��ԛ���r�nڥ٘�d�O�yhZ��E���I��K���\|eGQ�H(x��� �G-����C�Z3���֟��ܲ�2O�1�*d8@(�X!��V�j��~L�G� ��8LV����#�k[n�/�T��n��;�� 4�J�����-�d�����Ă�V�t�ƣ���VR6u��-�[l&�M5DՋ��ZР�U�:��&���$��B;�"G��f�|�7�j�\K��X�JMCͅ� L�~6~i"�}�L�b�a���S 8���%q:�꾁����+,;Gx�Jf/��^�vRū�s�%�zLMٳ�k�tU�xJ���g���lН"ф�f<J>ϗS�;��M��-�}�Dgiu���h	Տ���Y4�^j`ww�O0
l���}K�A�������xXu+W;�YO���	�%�NwY�)?�y9a����.�.�y�S,u3�M�����=���rF��r�uT��=�L97f7�� w���s�|����y�&���h��b�[�up�l�.&�ݼ����V�`��C$��1��ü�l�'µQ�i��K3�A��^^I�y�d/��K�J�E�I���iB�Q\����Aۜ94�ո�
�	�3���0IT�������,�O�B�QF�e�]gī�������'�K/����m/��`���Ke��+Q���i��i���!�5/�NC�#�!�L�p�%�`�Ӑ�]bǣ�v	(u��?u����m�%U�)�+UNY4P7?7^����?+���v�>�Ѣ��	����f���~��s����h�p�liyIm?�.�Q�v�`�҃�2��N�c��<�3�>9����i�2Ƿ�x�#̺�_U��\r4�sH;x_G�����]��A��]��������	�fH�r~��G������C�\ը�C��z�{�^j@�V���q�w�� ���o���<7����Z"��6e��ɬc@�B�f.<���,�?b�v2����2測u×Ze��Ф�M/b	�b`L8-�e�v_��d��`���o,�OF�8�����&��|-���0� �y��-��x2��E�]�7kCڔ��y��<|:�)��L$��E�jt�g�+�R�ܿRP�N?�mM8��0���(��ӱ`���V���Pj2?Q4��e�װ�I��p&Ɋ��WmG��p�@'oz��A(W�\�c������i)�ɬ�6��*!��.�,�~>���rIϜo�s�-�*W�
k�-���t��C�
��E��%f�F���l �ш�6����^:��jOS�`k��ͣ�1�:��V�T\��i��+}%)6'r��vl~��*�����5�*<A&�fc20���q �᫞]C�	�4��U�Ey�H�oT�Ӄ�L5�B*cg���P#�g�zVX���2u^����۰5�_%��U&�'�,�$��D�Nc���}}����+8����#��P�����4k̞W�3י�IiR�g*p��
*��`�cU�U��^��P���}��r��J4ۛC�5�k�n�ؓ�?4��~�&�6�o!Wd9�F��T�8�.,q$''����~N��@XÕ	��J��s/����C;��x���l�V����UY�ˮ.�t���aF�Ơ=ߒ�Og>��5��`Whhz�6��v=����o����
V�D�W����N�+"�+ŏ6ȵs��p��z�)�a���$���˃X��B���[��6��UM
��(|�����I���p�p*,l�w�Y	0Ǎ0%�\nH�h���~=(�I"ί��E8ߊ�UJo��|LP��xq�d�76|,}m�~{dV�<���J�غ�QC.��E���k$�jx9��yD�}I����j�:�dGk���@i�G��L�.�y��ֺ���=	j�y-�\���+D��3Jq�o��eN'�|��z��ܟ d!�G;�Lߺ�\2�M�K 7ڧF��s5��B����n��k}=�l��G�U�?,�#� qS0�e�$8�<;����3\�z����uv��З��³RWY��J�ٶt9c�JK���l�^'��#�Mqw�2bxi3�$nL9��T�_w9F�� ١a�q�}�����GJ���(E��0Z

Q}��!�$�(�!�0zw4�| �Q(3��W3�yp�V��Cr�c�iP&7���� Y��Ds�ˇ����(,�PH���k��Xm�?i�'ڪ�

��G`��A�F�0�W�څ�-Iܑ �h�xF�l6���	m�GO]�V�Bv�@E���g��PH�ZV��S�A\�����;�-xG4@W"����u�%���3���=�a�.=F1m�ϱ Һ��L	���ܘsZ���D.�T���q�G�d��"c�ᖇ��=�CM�C)�)���N/�*rZ�ы>/5�5Ш^�&�լ:]����]�;k+b�s $/�-+Q"z��}�-a	W�ˬ���iH�z8s:zg%J����9m�����A=Uz��R�f*�bY�vH�C���k�� �xR������.5x��)��K[\�!�d<~J�d�.|�P~�{��g����K�:	���#WMu1TA�=�@�hO�~��P� ���eu���hZ H�ݘøj����SФ���Z�\��b`q�X���#ۚ(��Zr����������T��9��P�E�\^�
&u�tk��S�6�{�YLw�yV����w-%�������7��A؈+�cb���u�:��Sܱ438}7w�f��z����^�m���{�C�!�>U�.%�u�-xM��4����U�>؄7�h�<�|�v�lp�?�f~*1�k� ¨�[���R+�4�)���8u3<#:� XZ��=�H��&�8����ؿ#��V)�$02��3S]�R�7�`^�tw~�IV?��s0bw��l7�1�������;M$Yx��(������r���MC�Wx�0��D�5R�%BP���u�WA}�隫vy=u���J�f(3ˎ$G��z��7*�ݛ5v����
\�3���B����dp��dK(�W?>��~zRgnӵ�R�,e
}\NAj��I8�+�k)�d�8)��={`��y�c��'��I�!����X��V��C������2h�f���q��ç"�0Eøϥ�+.y�v�e�h�#3|'7�=���.Ue�`*�;�O,���a��\)3p����5g��#�?�{�oS�%����wxW��1��ky���ف�'���r��$��`>@j�c)9RG̰E�F�d�d9��Rsk���L����ٌ�0W�f�w�J5͵)Nw+3&Z���p��[3�7_�-�1�|�(���]O��A!��܉�4b���J��VԮh�^���j�N��r㄁.o��jQ���p�zz|�A�rI��R<+��L�q���x���6O�ж~�5�)��Q��R
�F����&7�s��L�Ǽ%��d��ɵ�F�h<e���ܾ���L�ۊ��������^Ar	�:�<�1Yf��\��QI8a`�����% zz�}�U�5'�֝�3�br+�Nb��{����-a�W�	2�����w�_�?i��8;�}I�_�ܗ}5���b�8�Wp���}�cӿ���:�[�߁/���ܲ���Px�jS��3�+L�Rk]1��N���-��C)O�/�{�����d�S7t�	e1��E6;r�KB��O����km�E����y�&�����N�d��l�0���~"y8���?���k�4f��0`�z!@����8
L!���n`ki%.�t�]^�{�>��&V����e)�$~%�WL8¹��FWb���V�ل���^��u�q��p�fZ�**� �m�4���\u�i��͇��P�>z�^]R����:��v4F���4V$�L��<K]���8Wnm�v�GQc0o����?EMvu涼�l���{)q	*~C�E8<#�fN�^Ȳ���Y��FI���l:B³ ��/�`�1N �5�V�@F	�P�-��{2�7[Ao�x2F~ט�d@���	�[��tc[�=�f�k�XWN�QT-��=���ڲu�9�bZi��M��c�i��|�?����),���ղ����Q�t$�DI{�܏#;5�u��	~������:�$BHf<m�Δx��,�A'�i#j��R�4Sٺ߱��?f���%�ycix�h���]Fڡ��h4��u�ED5Q�n�� <	ql0�����H�3��A$^��-7?!�
����i��ݴC������4v��e���M!��J<70���WBc�{��;�l�r0!Y�( A���&z(RV���K8�t5o7h�5�=���ek��K���ZBq51td������UM�h�~g��c_2�o�l<� j�ܨ��?�'�2qz�1V�����1��a5���:��L�@�`�W���9r���ѡ�+��ܤ�����v+������B,�E#�3`�m�;=�뙒!�9�'�_��h�d�[��ǣ���?ũ�0��H��9#�}�*��K��i�G��+�>�@�y֖(WZ�Ms������%Bc2I�(שֲ]B�o�N���X�[���`�y׈=$s���J����v�1x
��"C��
��^u�0�;�B5�hmW|��[�>�������ZFdU˦�8��V������R�;G[�zy�,��4�oB�?��:�O4��^�F�e�g�L5�/��H�B���h7q,'yȳ��Jk��v[�&���&��$�[�@�~=~M�p �3L��QNx-�y��-�^D�������Cj���w�Y�jms�x�z�gi�u�*S�|����ȁ�&9���be!�O�Ѕ��S�F�jf���n~���(^�`*אdG=������u�.C 뿗��j�Z|��8>\�����<��b�����d��aɳG�Y��߽$�&'k��r���}��d�-03"~��$,@���2���`�_<S@"K-����G-�	I�1���b�9a���8N�L�儈�z�o�I�c�0�s���ջ �n*�SI̔>nv}sm%���Q�z�������5�~�^;�^>8���v�&]����e�$������L6vS����G|ŋ.�24��[���P�7�_L+z9���x��X���w�K���_0*�H !�^��$��]�	�e	��`�g�P�@Mu�Â�W j.�d3E(�!�_��
푊��RI5��+u�Դ�f�B'��l��[��w�A��r��=$uYr�:�tK=��qqg��V),*D��(�RT�Ƈ%�h��)�欭[�Z����iJ#����u
�!�Z^/�����~�T<n8���J��I&]^�n�WjG�����@�`G�;Ƙ��׋Ø���ݮ�u9Ǘ0!7����!8�Q9� cd�\��?'��g��S��S8W�@K�&Mp�~�c�qҀ^��	�
[��� ��&�٦=ٱ{�&��8�����4K��.�h��Q�/��-;�mY�YpL4�\�7��'�,_��y0 ����{ �y,�3v�9�)��ts�E�%j)n��DUc�����CR`��j��Ի�p8v�)@�A�A��9v!���v���X�O��B�������c0�ԃ��}^�d�l�����V	J.Q�.�e[*G�h�LC��>j�x�:O��Р� ��U��'�A^m��f�(�4� �NK�^�m37�CӁ�����8�eD��#٫�P� � �;�o��0�`���[�,>���n�.m̗)�&*��Ίk[�z�p�FQ+m�p�t-X�:�3�ɻ��f{�0j������՞�\"��|���$���I<�kkw��Y���+�~�3q.�c�Sa���_h����<��Y|�4�酻�S�፜�YM�/�A���-U#���QqD�F��2�e	��P_![���F%�<
�Tߟ[�UVJ��}���W` x��I�mP�m�Lf�NP���+�;:	3t �v��Ư#�XD}�����x*��k6?�QpR�=cI������M�#��>���TOz�h�]t�(�$�DS�����k.����Q	.��%�O��h}�g��\uo�.l�8�!�}rPm����rf�':�>%5bl�4G��Ǳ�;�\*4~R��*�jN���s���f_Ku������l��Р;]�f]:Kd^ɷ^	e�!=p(&�Lլ��q4e�􀕴�6�賥H� ��Ͱ:���][��>v7��:�J�2�b56+��KY��sd[����f+��Rs�Iå���Ϳ�3T&�	���ϗ��q6�hl���<^{�a-�YKG-���X6h�M�ܵ2��v�~�wa�3B_�J�x���s�G���*�N������yP�@QyO�$��S�)�X�7k;��� �i�5�_8ۅ�,"1����o0m���z̔@a<c���=M>��|o�� {SD��� ��)x���[�ɑ~�dn��c��G���� i[��G������E-ǒ���'b�h��Z$�9"�4a�^U���{ v����R�Ρ@ �0�x�=���i;�K}�ؖ�Qn1�	�1p�]����S<��A%uD�� ��bO�J�\���F6O�5�r}#��˰���᜕A�(�Ծ�5����0Q,�� \�L<V��֏1���}���WT����h�JC�!���۠�k�{(��^xc�qB@j ?�D�@.��r�P�,�NB�����ŴxӚ��L��m7E�n�ğw�$����y�9ސL���+AH)(<�������3��
״�����_n
�H@�5!cΌ��i�-�S������5��vDY���xV	��Y��i(��ZG��h=?a��:d��h�G�(� Jy\���4�@e�`YzͿr|h���.��^�gmFf�h���G��\;]GiK��҂��Q}���Ð|6 �F��6����<v�5�O�Sd3�x��M���Ols��dp����Ajt�U�^b
G��g��t�\�H:�Gw�]�\`z�}�+p2��&6��e���|se��6�j*c��ף�t����Aԃ>���t�
�f���iǀ|�In���A�.��pN�w��m�@����x札B�4���S�1�F�K
�>�A'mTi��������@X��K�댖�:�kb{r�	\ڃ$nMV�.�LTN���]F,�|����4������0�-�^�2�؆BcB�G��ޔ�����nm���CHb�)�v"�Ch:�U@��&��NŖ�'Y�g�?�l6�A;�1>1�qS7e�"וa���U@eE%��N3�6~��0��S��;wҍv�^H�q�kr�d_b>=�<�#^�&����!�?��sa�쉣i ���������ݧF&l\�nn�,n.C� ���*�����y��DV��:� Ѽ'��i\L���S2#��P��K �sr�e"�駩 �����շ�����(<r�%������ȩ�^������P���w����❵I�QH?S�����^����=wl����.0����	��5��(���M����3�J�ۼ��|j���S]��t�MV� g�VW��s��4�vh�q*tg3��i1�%������2�DW�l�z����d��Y����7OE<��B,�d�k��ΒZ�.�(���gC�o<�Fd_W�6����q2�y����n�!d\����5Q���l>9��<�a��a�Q��o��:��Tp��W�%<r�9S�x7�o���kU���8$�.�7::8*=zڂu���W�מ9��t�w��7ׇ|&�Y��_�L&hC���Ҷ�u���	2���

:N���(ѐ��hb$L�_'��Y�:\�!!f#���m˾��}�L�n]���ת}H �Cy��T�.k��������1F�a]%F�s~ �����E��:�%�gb�:ۅ��Ow
s�
�ܗ�l7�5TZ�$�sY�6cj�a��L�IIs�Of歀1Y���}$E��f�(1&���;�-YWWڏG�]jSkt�K��[ʙ'�M���g�����JsP"�j�B@w"�5C6�K�ߣUY���ٵ���(�Q]���t�ŗ��F�z�m|>�j����ko�V�)���$��7
8᪫\�ޫrM��pI�dvW!���X��4���������r�C������n�xê�f�V�����i�Z*�ϧǓ&�T������h��[��^�,���!d��&�(�yv������9����#���AP��`}�C��ՊP=-c�`���Z�o���Ua�p�1f3�<�-�aD**��\I�Df�S�!,��+�J:>�Qy���Rc��H������W�2��>1�ʙ�%J�����Jq���eM��
����M<�܈
�5���~g�-&�MH3�+�Y���%m���{���H�3 i��k7���b��(r�,� %γŀ���mb�(\��;�ݢ*vK#��hę������X_J��g���e;/3{�d>�����n�"�����l����<����۠�o���,A*���T�^q$��E��1�=0��!u��ꂞ��-��E��_�F�&�OWA�Pwc1�HT(�օ����������0�����VB�뺑�gM��5$FwIua���3Ra�������>�M��,�Jv: ������/���P���;��5�K����ګ�K��F�P�U�/�-�(��(��sN�w1�EO�(gǈH܃դ�� O��)�s������|���GK�.��3.��]�;Y��b2��cH�f�h𥜞���/�ܠ���`^�8v�3[	��+���m_�.�k"��n�+��L�=`]T_pj��^�v��;ٺX�I��Do�K��áV �QI�&�:��5ڙ*R|�y�~;�`rx)���TXbBGwC@%���g���|6�K��+i0f����P%�ٔf�E%g;���& ��U� |9l���7e�*m!���`$��p(�Aۭ��AJ-޵�R��J.����\(#�ѦtH�loD�I��
wA�͈�6,��
ⒸǊa���/& \N�X�cL�>UH5�̻�� ��~��0|���m�C�P�ضDYZֶ��+V�Cܟx��D��k���I	b}oW_{��0K�rr�

6ȵ�K1���|2+�i�������"$�5�[�����+͏�n��{����Řk��2�N��v���I7�L��ۄ�V��C�CV���**�>m|o���OL�vf6"���(��W����L�������čW���$U�.m�����=&4f���3cQ�?7)���n��l;��a���$%�p��OHk��l�aKD�O�~�'�څ�6�82E~*�"�}�)H 3����d�{��t�F�m� XVA���4)���Z��aF��3:<��l֯X��c���IZ���Dyb�C|R�[WkRl�u=��Oo��\�#����
۰Y�g��i��s��J���p�J�(�9{r�ē�z<>c\?�@s�r��W/j�JM��́�k8��b��ZG�<�\�Q>,.,2Q��������;��\�����vac�!}CK��W @�sw�2���f�M)��+	}	&��Q��+�{5��
���kF`v��h��Y����>�V�^�k'V~�.$���wI���7�ą	�m#�����"���υZ"B�T���)&
���E`D+T�F��U��_�TC�*��;��4�wYE�ZT���3ƅ�8���'�c��ͤ�C#�����./��R����y�h��d�ɀ4�4���^W�"H��$������wᢠFI��H\�ĳ�.b�V��W��-���p��u����Y��r矻�;L�Te�Cݞ�b�S^�m| ���=��y�cZ(2�*��T���AH��^։ONF''32%*��x����qu�e�T�=s����2֣B�ҡ<��]^���K�Z��|A�g�����J��"�D�3��瞝"�y�.�T?���)1L1��$]AY��g����v�����u`��Q�C���\���v�y��9���B�eaKAy�tlοJr죌�mPj�!V���D;��i���?(r���T��^�Ơ�n���1�mv�+'���\j��w�RWvѨ�A�5��T��qY,�z��}!t:X-.��(�hI܄�	t.��	 'g�v��ĝ�1�A�Y0���bdIܰ��3�VU�=�l�)&�@_!vm�Ҋ��P4<�4Ӎ6Y���va�����Q�qxuS��Z��M��39
���W�!��Rzn�R�?�\����x�1(�����ȭ��7�iky=_��T	�T�f]A�:��a��aֵ�U��H^
�}S_�x%�\���2�z��P�5l����G�\O��%<�Yq�u����7[i���$�����H�ɺ�1ɬs��X�{Ѷ})9x9�+8do�a�m�X�,d�:1��Հ�|�6vJp���x=y�-�.��ꑦ������:�����d���������&fb �����z(|O0�;����o�ZF��{���@�z<F��h;<���cZ�_���{\y|��~ɏ�s�g���>�C��R���v���{zٶ�栏���h��m�=�&O��!� !���+����v��N+c:,^H��e���:<N��[5��Ptn�^�?��I��坣���D�;��[βI��2�E]Տ�F1�}2Ȓ�^�8�ђ�-�i�B^�!������`�	s�'Ӣ�K�Q�×BV�	��	���ŧ��"��Mk��O}�K�厳�塬D��}q����0�Ώ�T �7��m��-��fc5�LP)r��2� #/�o���j����"n��3�.CTU{���0��o��M݋W Q��!cb������b��HM6������"�/�9�K��"U�>�t�����UoG �0�����f6]1"��`X�j ����4�	�|���Z3\�ᑦi�# [�xA�	��
����}Wt���B����5Hp�Z���HY[oℱJ�m��V/�w���Ok���[_z���p�W
�X�v<`�$۩��$��Y�q���@�$䔯����.M����
�4M��;�*8Z-M�	���h*��� �����&IӾPpG68@��|P��<���1����_]l��W��g<7IU
fsS���j�|�L	�M����q�~�&�u�������m@�ve�u��Y��^��H�K�M�,�2���ր�u��2 ���V�L4�9L� e�(�pBHfe����i�3��Q���Y��n<E �Bu���b���-U�Ga7!��רG��%<�,�w�5]���.�#@���[���=v�:�� nC�3�8b� ,=��x�C!�1�ڜ������D�A�_Q0��E�� HY��x$U,�)��8:�_��޷T��pфFm��*��e�����V�T���ɺ��b���n/�՟
1�Р�&M;Ɑq�i�؋�#n7���� ŕ��l�vż�$�\�~ju~m�G�����_�-h���6��N��(^��.�va�l%��ZN<<$�:+a%/�@��e1�;�����Dġ�F�kes�Jo���64衙T�sYǼFl��5�=�Cj6o���Q3���8fV�N���^ VE�3��↬(�sU��չ�o�����q)=y��ʷ�J�����vO���q��J�u!����Mؖ�1;AՂl�
ۗ�:�DR����񺽷��9	�\�����ȅ���D����r��X(�;�Z�;���إ�h��8�IRXg^"�Y)ۨ����?��Gu����k{��?7�m۝.)uǾ:�`�=U`*q���)�j�J��?_��2�	��6=]�pJl�5�&�jW)xў���ma�S��X]���v����I�<�
J~'��T|mЅ>2ir7\Y=G�6Dn�([m���鳆���
�50At�׫�'��G;��*Y��<�6������v�z�_觩/ ��`B#��p���:ނ�7���>��T�Q���Э��, n�sd/b^�^֤�V?ݧ���D"�{�A��`
���$uJ腼j����)�3j%.W�Z�HI���!pȚW�fw�3r�?�G4͈���e�6®�dӗ�t�
�ψ	m����6��w�;������^��p��
���]_h:������#G��oѲ�(X`��^�?��\V�zd���X+�����5M8�����9aq̝�]��@��f��Q��)�	k�e�����R��Q�@\08��b� ��6��3O��m�����;�S��F�UѲ��e���Զ�n�~��o��H���0���f��G�n��ma���>� �����+�Qw��m9<S$����U� �٧�5Pg��$�	�L�G����G�E¤ ��
�37�E�ڶi�)qX��
shM�?C~�v@����|s�N�#�A���D禦�6k�-�fT�dT�^��C�B����۟��ͪ/���fu�k��R�UOM���s#� �Y�� ��;8��#A{�;361�3��ϖ�i&� ��;��7O�i\�61��tL�q7�!��Hf(���(��ƃ�2�4�H���OЎ:��(j��[�雺.$�|]��r�iG��_�/�5=�|�<�_lt/��7�m+�_`�]681�钃y���9�����؁;�ڠ�"r�d��uJd���؀武,qn�L�\�SsE/��hy��Q��/���]�wդ%b4���e��??����<���?��%H���]+~����p�Ƀ���ԁL�\�\I�ɺ� +�7[�k����̄_mr�v�+���xG=��%ᄋ瞒Dhn����r�5�͹r��ϐuY���P�64-[l�� �,���Dc�B�3��@���)��Q�6�J�m����G;�=4��HO)��h���7o;��̦Á?DW�U��$��*��=_;�~�'��_��Kxnԁӷ���͔C[^�/r顟��ݷ!�^���l�l����`4��\^���K#�~��偑�uydMN/��+	Nc�D�(=&JI�&��D��u��d�!cv�#K�77MM�	�g9��	p	a�R-L��w���ǎ�|����()+O�3�����$�.�~4^�0�m`�IV#�e��7��Ic�@�5O��F���&��.!i	��X�8N�����]>��\�OJ��=���&w�^����i���n{xU>hY�j�c��k$Ք;	�;�r�߆Yg��*�&��<����m۶�R�M;�	/�th��'�h0��R���ދ.[X���lyʤN(x�PU�k۫�+���Fd�?��GM��{�hc>��c����У�ɸޯR��:��hS��h^�tK}��Zk�	we�r�y\Z�M����w�b9[ukN&_Q⽙�di����+���#�-������K���`f�;D�ů"�)ȬV�0�>k5'd��A����jcy�,|q��)!� Ҽ�$��	��q2b�¿>KR[y����z��%T�v ��B�}��-X�hھ�*E�B������_0�ʌȋ�7�5��p�i��0�����o^��߰4ҹ��*�y���l�_$'V݄��}Ճ��pj��e߯�i  ��5^�-y�h4{!�M��x�P���?OԔaA������RC�D1�h���~Y��3�]AAx�A�k�g���pg�Ahsb����v�㫙��0=`�լ�)&cԠ
l���"��K,�F��n��2mHC�j}g�u���d��4sʮ2��=y%���\5����q!d����.�}27�΅�p0y��� 3w�'��FE��\�ua��C���6�sB�b�q�<��U��H��.�=pAh[X��	}��E����=N�@�g)*����Z���w�V���΅	��)�9q`M�}��j�r��eQh�v3}�M�"�0N�>�h���W
h�:|�A�/�]N��<��<��t�
�F�OS�&���~��jO�iW���%�Y�){g���B(kB�{������́ȋ��3&*LW��Vk]۪��FB����;�]�F;��H����ᣡ.�;[	?����kM|��ɑ��^��;ܞ�p�qHk�%���zl�a2ӥ�X�7���m�HU��ҧ���t��u|�پTM��i��{�����u9���Pd��r�W�e&�	Vq��?��Mf `�H�5.6FI�E�f^ƚ}���p�_d��eL*�^��C������t���7;��y����$X'�Pq��GwZ�i�(��m���<:?���WU������R?�W!D��%;��V�5x*�S)�u�]X��_�L���2e.���y���E�2N���AKZ�mH� 2�/ �[^���q�k�X�A*Q����>��H�:Vf-����{[��r�1�̜���̶}e��Ro�����Cv��W�|��J3�>+k��HO�U�� ������a�'=�mK��SZ!!,�
�Ƥݯ���)⺡1@���vfZ5Fػ�/�w=�2s�\OZ�'��w!�3�i����#A��u��(�a����I�J�_�q��Mǽg,Tr��ǘu����.ď/A]��M� r��6K,c�5��Wn�r^�7cX$��@O7F(m������wC�m\�A�n��
[�y���_k��.�R>>WH5{�%9�۶��5h/ ]�ݫ��#�e �G(���8)f�9;r���g�O`~�=ר��!��%�/�
�~��ϲh&�"P���w���U�� M��#�|��Tр���y;�"�IL��B�?朸�^0Y�����.2Px�$ ~oI]X:Qf8�ޏ�_�x�э3�1� ���%��UЎ{�
��6�_�ʢq�J_� ��ǩ�?��n��EC�T ���iU���)�P��s>;f�����a$�)�JW�Ԭ"IXڱ(Q�&��<�ZZ��K:�O5}�#�V�@� <�Ӯ�w���K4���k@8� ��o�>��е�Y���;�#�LI� �1�Q:U���WOx��*u��()�i��GnV���� ���ګ����=th��`g�&��!�t�W���3'������o�;+A���`̧86�M!&4lv�����4U�Ѐi�d���5(��MaUa����j[�������^)�A�	���Z���A	Y��$����%4��U�� ��9:1�S�I�
��U��|w��u�x}ظ�*ɬ���B�V�(wf��cM-V�~5���U39��l�<�*:�aA.&��SZG������Q>֒�ft�	���]����,ڧy�UR����G��U�iV�Dlu�!}}��K���ߙg}������no�Q���AX���I�S�x{��0����CxrG}��Y�a/�al����l-;(m�D�zS���0;w%T�����*�����[%��RǾ�P%A#��.&�05�b$L<6�-ѣ�%E�UY�J�A���r��$xX�];A��WR�؁QX��bG\����N�o绌�("t�*N�(]��/R5�Q������=���3�b���HL��˴[%�TH�Gi�W(�۷Ba�o{��+*+:��00��e�CN��T��p_��< ��ąw�F9�1�e=�&��AoD����7J8����,�/я=W�0{^m�2�=���-��h�Cb���#BE �[����]��4(���Z�����-�u�~1���(y��C�H/*�G��!%+# ֱ�m3���f�D�~
C��h�[I�b�=r���ڱՏ{��f|:rQy�%�k*HAٿ!����v�J���$;�����X���%�*9�XV��&M��WE�	弥�hT.��8�=���K}{�KZmy�b�0�X����[�0�lg��n*z�ӌ7�f������ŷSp��Z��:�W*�Mh���:�xX���J�I"�먔���De��@M,��W^"BJ}s�� ��F��ր)�Z%����Z=��ں�]�.Z�D���<b���u��.�$���ilHw���-��K��RIM�����Y��~2_�/hwx#v�Wgd��b2�6�E�����&8��(#�Ȓ����o����fW�uW���^�a��b�4P�8�����-�4�{���}��h_��d8���1�wY�tG�ͫ��b���]�C�8�����D0��T���p�v���\@{�3��T]Ҷ�"��A��[�}�����w���d=^�؄Q�6�Y��,�`Q��5�-�C!�һ/�+����ͣ��!{%�b:n�d�� | � A�8H\���\�-���JUtl0)
�� �=�>�'�vl�ͻ�[�1�oS�o�Gdu�>oY� o�fǅC>'�\8.^��)¹j�	��~gSH�a�>7�����P[��4'm#��K�"ϳV�u�a���Y�R@���$�yA�qx�AF��T%�J�3;`n�Ys�����%vo y��v{d1�8�� ��C9�eS.m�J�,����IY��p�6��B7Fd�X'��ݻ�<ſ�x_�G���Q�R���La����A`�.7�\b艌��M�b}%Θ�~Y*��i!	
x��FX쟜z��謢�Q�e�1�S��
R8�9�(v���6�N"G>��}jCt�`y>�[�Գ�h������0y�\�C�;�����":���hV�y��,�R�GsR�ڒ�4�c�e��+"n�7OE�d+���T���KQ�.ڰ�i�~��<����L�9�Ǳ0q��?�t�)>��m����K���������o�4_U�������2A��,Ab�:��>p���ّ�R�=b����y�N�����Ig��$�>Sq�U-��]P�*4��JR�%JWn��bY���C`g���bMtzU�W��O%���h�9�Ҹ��o�V6����K%�5lݘ�����D�K�%P��y��(u}c/}9(�Xj ya��	��my�̄�GQ�����^�x%���(vC��Zg�������Lt��T�3|�Ӻ2���e(/1�E���0���1���.�a6�H����a.�ㅻ��wX �b�
M�U�T��p�rq,&+�3p�,5h��c.�$ZM��_d��C�%k��2�z�œ�Ɉ�sک��2����@Fb�)r�M��(oݮ���ȫw��O^�XD 6K�β�V��t �$"�V
��XXn4@��g�ʡpX��+�vݑ� `)����.j hCvVF�A����w�$��'DgRA�x68���Fӛ�U�EIu���������0��~��Ƽ�H����ض�}��b�zX�ֵ�V�T	$e��W:�M͠��XYb����8�B�%E����\�0a��Q��F�e$��u���	�/��O0�J-�Yn�7�р�Q�I�|Ac+�\ט�E/�4~L��5xL���~�iC?}F#��
*�v� ���1���<G�W�y*��r���T������ﬖ�`�壘�l� �F�,9�A����	�j�-�V"��(UZ-UL{�+��6�?�+'�L���=[���4�� t�j�m~;�cT�_p�ES۞5Vܲ�dl�a����(���w��"��T�*#@My{�����/?C�a��g��{|� i死6��d��+	O�v%�ܜ�$G>2Ӵ�6Ňx�\��¡!KW��ŷ�[�h�e�,�~�3�߭�N�M��`�-�qVL_N�[�p���6<I��)lτ'��c��6/PI���r�]����4c�w2�ڜm�Wq2�7_�֚/�%��
x���UOrY�#��Ϩ[�{,wnKp�Kq�[%Å�ɮ�ٜ$=��2h�-�"x��1�Mv��&9BlI��Yj	��x��=:�w��ʍ��mR]J�;�#N��j�?��ȇӁ6b?E��G��i�"q�T����1r}�x�b�ρ2T�6]��a涴����,m��D���P��$5l���8I�g�>"/�=��<���Acl�!�m)�`a�\yc.��!,`�[๪
�.Sq3��� �)I!vQ�b�`�����`��rЮMS�f�Q[Ə�b����*�r,������~��9�)�L�G����w��ȹA7�9�i��ʁ?*�p�*SN���a<P��y�3i]Q���s?T���5�Pb�B��蚦Xb#�pv��V	��PejqNe������ָxϙ�&���=�қ8@�3����Kiw� UNE�ڽ۳Ue�ן��W�Q(���7q�G�ka�S���Ȥ\)����L�($��,�b��>p(|�N�15�Ĥ���/�]��[��#�E�Ft�����He8%`=�G˾Ԧ� S4�&AgڭO-�ey�j�L,��ٸI�v|}�~*Y�T!�{Л�[�9�xg:Ü��Y�����ӈ��p�!鯞!�)VQEJ�W�c��0�E���J��e!8Oqe�����|$]��l�7xBX�İd��XT�QgO�,�{p�>/�%e������EZl@���.7�8�Rn�w�m+pT�0p_7X�X�<�)�6Њ?9��I08j"�[X�CW�8;�������эZ�8�!,˼����p��a�F��{-w�*OG�D�-��W��Ӷ����v3&�5�r�}k4�p�S��;�@�(�K䢪���%�r����|���-X�s.�����R��1�R�9�ΐ�dwN9���JUF)u\*"���yEE8�W���#��4����~|�+��Nl�<����n�N���&x[�q�Z���1*��=�������>��)�������&�9]z��L�w�!�վ���F�x ��%+�LPA/?��5����3��Y�s�w{XJ���wwp厈��l�A|Ҫ�=�c�7W�����^���Aq6��o- ��y(��� ܕ_�z{���=J�,KK�N&[5#�1w��KO�tՒ�N�p��]F�C����!v���Q��H���މ?іmٌ���BY~6V��װof,=�����x<�EƔ�$��dá��@'���Eyr�t,x�
��J�� &T+:�y��,��nP't%���*���7A�=�	#j�x^�/�$o��\�Yk<]�r������u��3d�o�gDa����se~���r����B�st���*�GI��0
�:�Ʃ��h+o3��D}��E��^"W	��#��+|��A���C��e
��I�;������.���Kx����!2�L��M�RW4	�߾�/ā��X�t���<�o��x�U�|>�M�z��7��O�q��T2��~���LI2z'f ��gwA�?E�+	�@+�Kɀ�,��Z��u�w�����j�� ��jc���Y��F�,�N".%�.�XP������YYo@�@!�0�c`՗���"ue$<W#0@�ܭG���mY����涨,�]�֠,��l��\�a���6�T�|˔��9R�)�/(�dC�
dh�E��tj��Dr2{\�v�q�����Mk��:�ܰ�&-�m�F���N�2��g��ٓ����> 
�dLA�I�XIΫ�~�m;���
�N+o��
i���0.��Q�"�6���
������[�����K]GO��������r:yBH�u�@&�r�0�h�;L��3z��Q��6���ӁK�=���Uk�3�v�z�s	�˘�ݓ�\������1nYƯy9
��=v&���G8Ȟ�{k���Wuf��ď_��i�c{O��̤\m�5Te>l$T��i2]�@˲|����	�S�l؛)����nk�?�Nk$�lJ��5���B�$IV��#�DՇ�����.�v�O�x��Yz~o~p��IUA�V�P���{l�M'oN�
G�����8[�5dz<����`�3��7����OQ0]���Ihrs�E�g�����_�����/�I�Ƕ��_Q���N#:?�@s�L�{Z\��N�X�	�B_��2���9F�C���*�ۢ�8,�	0D�;pY���e^��}/-`�;���wj<���3Aj±C��j�����=��Cx��I�E�̄���qUD�WK���O�"���hcpRVt��1��HzGxW�FyJc��C��E��Mh��ԎE�ڞ,��aD�%�����^�
%(G�0��0"�>`L��A �O꣙��dN�A�SP�$�ߴ�8]�����fWv���J6L߻cJQ��{8	����o����yIp��!���,�+Ki�4�@Ę�R*"-��D�����
�W�=����QE�G����8�Q^�pH��xN�I�}̦�3]g�(����i #�"9�������,����Vc���p	��ph�y��-ݳ�..�.���l'����BBq1y�Qe񃺥Y��7��Dj̥�}ªf��tz֎���J�=��V�@.)�v$.R��U�8;���KI�<��p�����1ӕ��E�W��a�i��Qs�`�n-�H�/O�M�n,���� �����A�xU,�Q/G9�!������R���c��{��J������[����|�=�|Q�"�C_��pN s1)3�i�h�/@�f3��r��U�~�������g	������P�q�m�O �pu3�j���F<�d�������M(z���N��	�ȝ$����ݴ���U�ם��(�=t���_ pS�"�]�ı�?(Y)�T��QF���&�L}s=����j!�(��-���V�r�+wu"��LO�w�7E����A��Dz��S*�I��Tۙ;����-i�"ɰX�֏49��oq��NR�0,`�ރN�r��J��@���d�"O��m���Ry��]fb�6���� ��"��y�~��ёF�1���uG�e��0'qq6D1G�m�7xr�\)Qj���ޮ�s�mX���벿,;���<���B,N�(#@/�L�82��h������<�k�._�9�Gp�u���k��?�����X�+^���Wk����O����'?�p� �����
ɌE��!Δ
f���p��k� �
�A�tU�6o��|8ٻ�[e&��v�=˴+�h��#G�����U���I	�j���F:tsf�ȃk3Y#<Иc��
Iّ5���ƌF>���tK��Y�:Ov� \���Ru��D�:�.�A}�*��r:�b�.����D�2�3��{c�Z��&��@�Sr�����*��m�v��0�m�1�m^�\q��Bb-�
�r!Ǭ�b�f�.s�-g�3��+&m叁�Ct��T�DC��d�x�[>�����:d�c��L���`�1�GKw81�����N5�$/�5-F��E��\�iO^,��ƺ��Y��#�����;"��Y�e৞|r�T��%H�@"Z���s�����҃�.���5B(����G]څŏ���w�A}���>(�i�\�{ѻ�����(�ߢ�˛_?!_)����P3�妸 E�C�7��I�~2�s���t�iU���%	%y�p���:Xi��Ѣ��	����u��-*�	6�#9���b����?UZ�#@�g�C"J��?���=��:�w��+��_0#�~Џg
(�cL?F_F��F��4����1��h� ��/��?DIA�&z�i(���_'t�m{��:=�S���L��eu� ��-�("������2GS�$����w�à/�GV|��䛟�2=�����)w=��ޱ7�!����[�����c��(6|!�;�7]zC5����q���J��J.-�^��|�6q؏��3�׺k�2A2N�����B|#�P�;�+$��"íi&����|�k+�Ȭhf�x=�u�R��L��ǅ_|����)��B� ʳM�ס̒���@��^_���]4��^2��Oiu ]�!q���ٯ��g�����c�S��Og��e�fjV�����=5�MyG��¿3^Tn��\T�O�,B�M�(���٦L����Hwt�*H�7���ui��.]Og4!����M_Wc2��Y}��1��pQ����F^w!v.��$��{NB[;�|��ps���ևz���J�6pn��k�)�i��8wX��{R��>S~юz��Q����*��w�������k�#�6Dn����Cq��<�Y��>tDx�kTr^��lA�+4럼�^�j!�_+�:��!�M1�9�vVeNo���K���S�a��H�H�2�=�t��|F�-���� ��8D�祋���	.�{5D��&&ag(=R )���w�݆F����?s������O�H�w!�vf>�dէ�� ��^��~��ѼF:M,�p;�����:I��X�p�n�z����窘�ӹ�B����}v5A�sr��	* ?1|"��v�����eД��)��ִ�Z��'��
��T��M������s�)Gw:1�$c�o�� �VMuMi�o}l���'G���AQi�>�g�=�����8�Ov4�JZ+ۥ��yw~�=��|b�]&���}��мH�5ڴ���^_5�����Y�*vS�{�(�ǒ�\8\H�b��V�,4ݩ���t|�=�	��|;�ix仜����j}m��~�'-�9h�����������[�-Bo�%�x�O����'�*I�et�g���G%zˮ�j�Oظ���T�d�$�s��ss�w~�ZV7&��iJez����i�?�~���^�*��Ä�\@��e��$�&���L5:�ʈ�s��7w�V���7X���E0�T���
|s�����޼��}��C� 5mE�m	�y��K-o�ǲK�	}��~E �'��mp�σq��w�j��[zqk��Z��6���Ҹ�)rZ�O�7h��C�e�K����N��O5Pb��-7V}fi�iྀ��}��ȧ'MeTR��霌j^�a/ٴ�������S���B"�V���b����`G�z�Ɠ{Ga.2?�l���kλPg;���qV�R�9�q�3"㛍"	���f�i8v�~������Q��9[XQf����l�� S�z��E?��Iܰ���Ib~��]G6r�	|�M�	�nGc�Rc��܏��)�--%@�wӺ-!Ϯ]�h4[+��I7����=o��=��:O�%�S��;(c;B�<��\����܊���%[�}A�����ddvo�����t�哢~������h�H���Yǡ���â��1���QBʓ��p1��6�}�e.���7|0w
�����p�Ĉ�w��Q,q�&��H t���M}���Nm��;�u�f��H7�(��ALc+�y��[EU]1�3(�é{7� ��/�&����JN�c_!<����:'����!݌
��B�%��_K^�]����A����W��4BqO$թ����%�4v<;����7�����l����j`4Gl_8�ۗ9ؾ#��P�P'�$�i,��Z�em�vý�H�wb��� �`[ս��%������0S}Aw��Y��i�fRL8�Ε�������t�w=�`�Zj�����^�c���K~q�O�����
rΟ���p�I�1=�ۏy_��{n��
T���!�WD�5S��K��w�W6���o�z�����v����v����S�10	K����M&�H��zAQ��*1�\���.�	��(��-w)��&s�_x'H^����_3�T�����Q�fn���߿�ȡ����2Q>�������j��J�S[)�8$5B�hyvD0��H�ZԊ�
���	!z�?�e���맱-������u�LZ�EҾ��C����u`��[��D��P�)�J>i&ioB��q���7���<?�[p���N���?���W0o1X.б���$��g_��|�k�gt�)��SVE��P����6yZ"ָE���~So+A��K���Sab���	z�Io��:��V�������<aCe���8��p��m���U�y.4|7�0�z:Z���R�&'�|�a	?��ܛ:*������'��	���M�]g�Ȁ*5��:��φ+����Q�D�\֝���Y�g���%����ކ���J��䗴�i��j��$B` F:Z�� ]��U�%�P%�����Ԇ��L���o�nlY	���#�c:�v*)H��ay#�|G)E�<c�F�P�&��b?I��h�+�|+a��w���"+��$����M��Q�\N˛T��H�[X
�ޙ�J�4OY_�l�\���f$6�^��3DK��9=��4d��޻Z�D*d�875WB�&y�u�C���D�L�vuN��L�!���18�h�_�����5�W�J����پb?�>��͹�� �!a�/�v/��+]����c;_������S7�0h���v��T�)�B�I��.H=t~x14�[d�YK< .n��XH��-o,lHIX��Q��&#ph;I�p霣���䵢~:�(�CU(�{mE-bJ_#)��թܞg�攨�/�$����ᙽ�A��������`�����Ƚe�4���|���Hs�j�ѧ��mM�3���y��'=k�H�Ht�η�E��V 2X��~9v�i�DX�?X�J�A�r�E������+��n:���
γlz"2�JJ`���v��i����K˰y�>˦�9�s����jI�/ӱk}eZ�F8�Ð��K+t���1y��h����
���E�{���"��,���o�CӮ*�nM��v�2��L�O2)h�\�QE��e�n@x��(�� ��G]�k�An��M4� �z�P���T3gբX~+{�U�0�	��~�����v�>:N�?M���"�R/�X$�+15Gιa%]��Q��Y���LA�H�{��H�b�4X0��v��?H�a�0�2��O�{�N�q:2}�;�*3A��b7�c�,���>e>k렢P��O�φ��O��Cz�������:�����?x���~o���ZCֶ�Ø�f�!��_*D[��(�p��9��3Aa�<x�$JC���KO�����ˉF��|����C����iI�����Kp����j��?JpE�·^�o�=�m��`�� s,�ƿ,+� �)�p0��U�Ӱ�5�P��3Ī���@�ٝ��I��*f���J�JD���Q9-��L���,��ʇeK�?�FG��U]9-@����{�*]+/��s��d��t�T���baH���=U���P��3EqrY����"!�#��N:Z��|��_eÚ��j���-��D��ߒ�Gg���գB^�6�
7Z������Đo� ,�p���:�BuM��r	��*?��p�_�ZP���wD3�5d�y�3�����*��؇����l�"-L��ߝ���`�wo#���y��)����d��6��	:��k[����²�d��)�p��c+��ȇ[���h�,��f!���;N�#�{~M˒h���%o4PD�x6E-g2UzLZ�#�F�Ʊw��0I"�����V��/6(P�'&4�ύ#���I2qf�+(E���4�贪�xT>��G/�:�s[^��~.h��viB�z�870�#	��7�]
i�J�;_�QO[���nֳn�0�o����8JV^A��bO��w��5ba�.�y;��sVͺ��fK�?�n�f?�$X��6�@���&��eM����B�tya����OЊ�v�4�����V��Yz�ۃ�Ğ��v]�Bi��}H�ށȼ.H�W���%���Y���n�h���L"����� v\�~f����[5�y%��<��ĔA������p�/�/e �n��9�����|�lc��ꪮ}f'u�,���Ʃ����{��U����TG`&�S/=G/��a���f�_�0.c��M�lﰚW�t��N�f۱�oӕv���ʩ)�Е�͖IP�7�|��s��L��ΧS�
��H)?��̮B�Nba��PI{^� { A.�I�7~�>�����9N�.zء�q�A8�)Y70�n���ŰGo����M��d5h]q� j�F�#��w��y�2|l�=l��B�Q��ɖ����~����D���B=�[��s^��'��eM,Ü2�WS��a�J�	�Q��,⩿z!����)�8�,��
oO�K+ZV9&(���U�v�E����~��Q�+h��)Erkm����7Y��C�$�4�u0�0d��wh�V��hYBs�1�_�����E%�w�t��{J2�������5hu��X\�%Tc4j5��9�y��� i88	2���R&�?!H�|~���K���w�{����뛵�@�Os��@� `f��T�0熮��S�4����|�ߔ���k�0E��g�W� 
�1#h���`nN�
9Z��a4�2�F͋�ũ�c�����f��Z9�?�ʦ>��4K��k��	ɿ�����R��%�546�7����x�9�|�u���h2|J��j�U��{�ҸD�1�"�Y���-Vad��>��n�jLa@��վ�蕖!M�vȾV{R1�ၽ�ǉ,����W��:�Rw%򕉻��Qm�	�:]�Ʊ{\���-H��u�ahZ���T���yɻӃ.�l9�)y�0��KSN�&w�7Y�T�:�YfՋhN�3��I���G_��9��z��ض��r���I��>�����^����>��������]�M��Vo�GT$��X@�G֙�e�~6��<���%����#���Wo� ���HK'��i�9�j�8m�k~{��<������3�_���3��y�l䍸r�(/��C���ܼ^�_���Y�&�HA�3���ݲ������>o4]�g(Ͼ��!z���a�,������}�(Xm���ٍ�H���ۺE�@a#EJF���!T�m��TS8�P��0I'6c�]�贏����4�0}֢�^���S)�m4��T���C��~���s@ɍ�l(��3n�� �it��m����)Ϊ�\�$�n8�|G�V��* ��1�Py	�N(c�L��9�W��S�� �3��V$�r����f�Q�<�l�D6k�����ȫ��zg_c���H��c�5b�s�$�" y~�la�=Nt0j|+�=�U׏��xe{U�E|s���=����a@��uO��·�n�9����O �1v�������뽸�D��t#�� ���%�X+�e���;q��pe^"�pym��(]�I�ۙ�F�T�,��3qh�ZmR��t��JŅ�\}��|��uށ����O��Q��m:a2��Ȁn�0�8����rB=�����&-�P��9��nn�,�mF-?5 ���S�W��A,C��Rx���]Qc,BBJ��)���I&�c`%��G�����E�k�ɜμ�A�A�`��k$Q�� ����V�ʶ�<͍i����Ⲅ×��!/T�l6�������FP�9C���΋Ƅe���[�F7�KK��sf�Ôa�$�T�JM��^�ג-��2�1�#ä���'�2�%�ji���}Bl?��^��6/�ĝq�^{��(So�'Yzl�Ԇ$j��m�r�y�U�M����[�����ʏ-��U~A����#UBK_�p�'۹���������G��+Q�*�jo�V�4�mİd�N��"szm�sOHZ<ȁV&�ٛ�"I`W��&@[�6�/ѷep�n	*|F��w
����������7&���T� ��je6K;�'�������<�x �Iv����6��}[����smiiz�?�9Ε�i}��ZuI력7Y*�RK�_��H�k�l�*�Vi�B`�/R�1�8z/g���:F���^�������\�t�y�	���a��uݓ;
B��cv�◷����9�p��������"v�PO0�E���v�#`����s�P{�ƋoBi.�:�U��pzb;�ѻ.U��B8Mivd�6����	8�kf�d�h����O�W�s`�xU�7̑��1��R��S�Bz�M���f��6�܁G"1N��Іm�������n���!/W�P��_P+��H./,B���ED��R[8C���h?MQ/�4S�&ݬ��y(Pc�F+(]���K�iAr�tl�oz/���5_:I~1��x:�':躄���(`�Ӿ�c�T�����5[��j��w|u��Hp:�	=Ǉ+ L=���v}���iıL�1m�Ť/��e¤��rE���N�L���t��H�be�
�?ue�K� �%f��A�f�!��x���<�ܑ�8"�RͭδWrk�N�����$��d +��g�!�2�o�HR������{w�r�s����E��C4k��΅�6�n��s�B���9U�#W@�T����v	�b3� ����/�@�ެD:i��QVᤡw������
R��=~#C�s���D
�+��2v�����E��O��T�ie��É�n2�QZ(�U���潄PJb-�oa��8<����]92Ƶ���B��D����v��	��*��eRk� O;�_������3�(VɰCBTV=�Qj�0[��8���>���p�-�uR%�h�'dI��;=o�s�h�xu�{�w�;�ѝ�!��̋��vѮ�$��E"w�Y��#�ے��Z%��㟤��Ho���v>�pF��|,#2�X����i��j%�&���Kp���֨0G�՜��T��4���^�?#�!�2�zh�8F!��Y?F�E�����C�RUY^,;�s��� rT���ЛA�kn{ir��j��]����<U �~/�y��*][�����*S�Ri��tk�m�ݿ�"����RL!( tT�P:4�F<Փ�Qg�\(�\��cm����ftmw�aE"���f��;;�#�]Et\����nm�|}Jq������������ln��;t���/��<u����}YH����+��̩�b��Il�,��xA��KL��&��ɘ��5z�Z�d�X��-Y�Z6��S�+Rg�%e�`�j��O���u�Ʃ��u�����/K2.f�����jL�����b�gu}�))�l �pc�?���FEZ�Bt8���w'��%n�ˏ�;C�� uѣ�|^�?�V�F�����	��;��$ȥ-���˅Z�)Ff�x�PF���t/ŏlk}F;�o�@������1y�k�C�g�P�����ՙ���������<!$"�E���֪GZ/��S.��)���}�Z� ^F�B�􍗤�R�D�V.�ˡ����A�0���Kdr��݈��@P6	$5�[�Õ=�|rvO r��v�8��p�2s�<��-~��^�f�������όa㐬�{o*�L���0�P�Nf��/����o�ȻH7O�t1=}?��^mM�_���ee��@����~4����l�  FJ
#HT~@�
�]YQ�6zb�g?�t�`(퓬�|�i�H %#6�i��c\���Na/��zI:�`0��Ǚ/^e�_\�* �f�G:�?l���d�����q��M�Rcx��*}���f�*N���U��,��x��RL�&n|ҧ�)��M�u�`WO9>��z�Ȋrp�$��<dŅ��TD��?r��[_��W�I�G3�f|��>T�K����-ز9�rw�2�X��KL/J)�yͲݓ�J���lP@7�!��%[���_�^M����ř�.���5�f��Y�e�=�s��Apq䭾���_Q$������k� )�ݔ���eT/f'�iҫ�I$�ykr������ƴv9m�a����4�O,��<I�S�7�Z����H3\�A}"�9�č���t�&�5p�需���J��z.�fX
��[�S��G��0Կ���x84�^%�~>�ٕǬ����.ӹ^�D}���òA	�n`
U\?� ��d��,I�VX�ņ=aj�k`ɒ[���A�*��<`U[�4>�W��]�k�~ך y�W='s|j�B�ӷy��摵�����a6�C�6��� %{��K�����N��g��1n� �6�YN�]�}�7���TH�9E�&���JG�%M�|��p�Vdݓ-fs�L�o��z�02T�z�g��WU�/<���@g%�V��b��8o�Z<�3ܡT�*{]��ɘ,m��,���Y�5��"�nU�Qm0��h�ȭ��(A���A\��n����j�ߜ�������������̆�������HW���d��γ&Ӛ+���R�F|}A��;��(�?�;�}^���2�Y�������#�I�~��f��l�PdX�/�(�	?fJ����^
����X!5�/t̖�u�d��(P���o �����+�?1/�[�� W��ղ�1e�Fu�����拁��z~��Y���'j�ս�����6)5-N�E*d|�\�1���K� b:���s������4�~qy-�2�*��\���Ƒ�VYu�H��Y}ء���o�֐�$�B����K(���FR��� odq�G���e�w�m1P5�W>7� �a��r) �S�t�iPa�xb�0��Iwp��V��L��.X�i�$+��b���C�Hj���o�kA]5u.�H"���Z�~�('ll71Y!��衿�V�u8j=���/g��xg�^<�*qbF����R|-��f�y����lڼW���`x%��z):A���KhOމ��SǊ��L'T����N��|œuի�c�/`�N`\��R����� 콶Pw9�6
�=�u �m���5_!�⬎�.��XRf��w��r���.�#�hU�=1<I�����Vˆ9�?7�����m�+��8Pd�L����5Y�r@)�� ���Q.
���d��'�=�]bB�;�ԻIy�Rf��F�2_�1�C-�;��4���v�|7χ�<�	��s)��.58k]��\}ыd1i[O��LN<�(�R'}} ��&K�m!À&�|���QŃm4Ey#�L���1����7���*���:��%|���X����k��jƙݳ!���$��[��l�{�+\P�zE��+{�V�E8o'ěr��������!��Y�g�K�c�ď�Yx���)2�zZ���O��D_o��>N�S���|�@���
��^��i`�2ϑ,&�v5��]�֊=Cy�0�e��pةG�
G.BAt�IQ%v|Kg�
͖�H����*]��n����&2OU`���V��}!h�a�t��(Ş�*X��ȼ>}iU��"�w�ψ�}��tuL�nR����U�.�Q�2�Ν=�_ _�v�&J�s�0�%�]��S����Q�é"2����ײ�U�=M�#5�wa8��ewG��Q��Rmu�[^�^W/h6��l*i@���P��j\�_\*���x�\���ԏ dbf������4��8ֶJe'<ǁ�y��\Jna�ZH������;���71����4�r�E��嵀;ƱL��j�`�^Φ"�F~���祓��l�.�^�8����������;�7�q|�=X�����ȷ�}�����T�6��qՀ�ӗ2>�}=R�����������t��=�1r�3L��z�Q� Cm�(l̉���M#yC�ͮ��Q�r�������TM���K�B�Zn^�� �c��5�s>
 ��>!wI�q�G|���|�;˝�!c.5Q�T�y�̮7)��aJ�U,���21��3;� ��`�YɎ��_!��y[b=L�'�DXi�i��+\>b��ݨ����p��U�HzG���s̗�D�&�_��<	Y�]a��$lV��9��C�:�9nsc�Iw���S�R�w��WS��tQ��1o��������UO6��;nCЛ�@}�<q�	���T��@�ƛuɜ���O�%	�|�EKϟ�������n��i� <�Od�d��2� ��O�1�k+�7�_���]�eK�W�E�9kt��S��|9I@�}�+zR�,����1M���DQ�+G$n��L��3q�0z��*ͫ-侉X��	Rp폊�����)K�,��S	C��ۚzO�������Bx�/��K��<�#�Y�����۞�w�*
;}�@�����:�2[+55����|č���^����OiXքP�Xa�$[������&�I�b}!G����.6W��pr�8�ɜ�Z2��8�X�:�V�sx�<��V�����3n�4����s�.��o�i�@����2a:�7�|�����.���^�S7p&py��Q�'[�e1i�f��1����Ağ|V����Yi���W���={@5�X�뻣�3~0�j0�Z���KE�m�Dϡ����<ZY����v�MZ����Aq�o�_�d��p�p�?��
���L}zCZ���l�
v0
M�򪑏H�q�{v'�$7��&��(z���|qU�v(���0�'����%�hϼ�,����Tm�
+.���X/��I}�Ժ����Z�\��l���g�l����C�fk�o���a÷����'��Y�+�����1�(N9�H:磃c�Ĕ�p���*�9gy	��XQM|21Q:��X�}�wCT��J�,�v-I6GՂ-D�5夭%-�C���d I"7Օ���"c"F��L4�U�[�;�lr�����dJR=���4�^�,�w6���@�P�TfQ����j�ʷ �3(�:#sӧv�T�V���ﱼ���6桷����Ά-�ɬ��W>�9D@=i�a��?��u�8��a�Q���ۑh5Q��8��~}+\0&Ī;���� ��j��@Д�Qxq��32�A���k`�������R1Ǒ��կ|����@�ۆ�Ah^��p��Nkv���*��q���(!�m�g2-
��{��x,3d�A���o���E/Ti�i�p���F�̂�
o����{k/���qY�vD)�LV���Te�z���N7&*CO��y�ye��{���5+]m�<���@�U��Hؑf]� �\a��§.bn��u���`�u�N�����o��U��#B���G�e��Fg��o�/
5��d�ޅ��M^�t8�8�h��O�1�0xF�P9���a͵������7_��)e-�FR��=�J��0�V�]$7�* ��j�K�+�[��\P#�;e���J��@�0l��A���wi:.�������ݲ�I�̌7�NZܨ��G�4�3x�k���͙n��Md��-B���%<�������7N��1�:��p�59lTOgBNA��Me�\�j��}��"�o�%}] _PD0��-w���U)U��B�PsU'u���&h�z�x��%�V�*��F����V��}eqr~*bb�[�� I+���R^B��Dy��G$�0�C�*�WV�[^�d� �z^�$=����&����WT[a_
某d�ۗ"���Z���5\�L0�a9����m���b�9��,|�b��~�h�&�l{����h���	B}O�X؏�՗��21�7#�~�!��Z���=��h�����:#��c��M]ƞ��˲�u�K�ۤ�j}�US"a�$�,��LT[���7��GW'�����uV��V �������=�}^̘��J�M�'��|'��6�o��T:d2��wB7�+al���8�5[��KF�:�k)�3��!ܳ��B��>�t+'c�0\SZ83��B:ބ��@����h�d>e��p�	F��^|��3Ţ�f�ߍ�?�[�4Ͳ�P #y��2S�,�����qj����#vv�JTt�,�21�y��� g�E=�*A�q��:�v0�[�n ��]J�{��ԯB�sl� ei�T�0�`Y~j��N�Nv����O u�i�0e�Ї��#����vf�<��fمZo:7���P���&�inV�t-�牪L��Ҝ����#����1�ljIfL8��N��:��vRwݒY�"9����%���i�V*��2CN��A��˼		���8��(b2hJ�џ!�XC�$.d�<���G�^�H6��]�$�g-@�k_��&�E"�)\��{~io��h�H4A�L�ƫ�Dň\?ᩎ�{0r3(�B-�z/`l��U0-]o-0 �cW4��Ǽp��P� ��
V�˥Hk����)(Θ��뢅(�ʳ��C1���ؙ�[��9��O��8��Z�*����)sc�i��"�G���B�3U����9��ў��}����;�m��*
O��L���T������'�ʌnQ|�.c��+�ߢ
x��/�ẵ�&�4o��'�vi�f�k��pA�,,��ǫV�&x�$'$��^�`%^��_l�[6���Nރ�s=�s��xc���fٲ!��W�p����M����D�\?��
���N���{3��:B�xf#:]*I�ߩֽ����F�UD�ʞ���
�R�g�2>�~�3!ܢbq-����@ c6k6�%C,=Ń�; �F�M..�C�-��,��1+�axګ��T��Zĝ�L�:xP�d1�(���&xcr�I+4�������/GŞ�����!�(��=������i7|\S�`�L�iR)w��O�I�ͤhd^���2CW��� ^��l�q�6���8[�t�8�/� �
��!t������Y�znG����ʝ����<�O1|��/N�H�����ؽ����ӌ'�\��K��Ѹ�s����D�d�psek�7�����ҦJ��]KV��{s}�G=�τ�Ӛ���cǣ�<J�j� fD���<~��H(�����p�y}�
{��GŃ;7�Ĵ�"]�x֤b�6���c����7Њ�)>�/�<���,!y���
��4�	ߓFo4��M�	�z�2��j��|��(��D�1��Z�w�i8���}�&d����e����ɴ��|o��˳���C�l�����'o
kwFj���f�~M�r�
Ӡ2p�,�6R��ۃd�dB�~o���'����7r��%�6\M���s�H�:ﭭ{tڒE�h�'\]�h��gQ����ȓ&Q��h"=������[���?{^�0nD���6�',��I�
���m�J̯�r0�Hu�	�������k�Mx/P������3>����޾��d4����t�m�v]�Cڼ�RH�~P�(��f�ם	���D3�=��ۯ&}�'d�ƠUQMC�"bH��c��O�-���Ů-����@�vz�[�d���~�xR�%�����v�D���>U/ay�@[k�z,sO���� y0�Ƈ�t��u�����fvT����ۢ��9���H�����'#��*=/;�3��������׌%���u�A�'�?t�a��Aµ_�)�J-���&�T?($E)�������Ӂ���
���7FL���,����;��'�!*��n��p�8�3���4� ����j�}���`����8+�^7��4�Y��nr��zM<4ӄ��Y~�\��&�k�����t.��ӣj�5h����k��D�Ųj�����yE�?L�ϗ�z�p���?a$�!Lpڗ��n���gז8�I�;����r�Z6��|*��߄��P��xN[l�!��p��&H	M�W�K�1<�����U,�E%�m�(�����D��o���� m�]�B���e�(��)�F�?�=ՉSE�#�H��U�) ~N~ҹ�U�/��p����T>���,j�=N{xݎe$p%`ˡ��}h�cڛS�!C傻J��j�&K3�	T��z�k�%쑙��Rs 7�U�
kt�LF��"0y����ːP7NC�/z��~��`��9����hl�\��9��~��fH���ﴊ��|�#���Xj���\��(gR)���	�F��Ő��L�g��W4�5[���j,𘑙��Z�B���_R+,��Fx:p��)�h_��sJ�'J�R�>���'�ZY筋&�.H�w��oǽ�`�Xi����dm��_��j���n�&Y�c9�P<�d���wě�+!v��`Ⱥ�[E|Nel����V�>81�CPeSCC��ۯ�ɚ[/[��c��^,����ֆ_�ꗿ��V�y!��59������avt4��8�?SV`l�Ԅ���\�D�PC�qo.ܼ���B�q�29�������s}Jd ?���z{��S�$
�T\y������x���Ū�A�%�?$��g�N�Б`2yU���o���E����I�c񷘬�fJ|QϹ�o��}�P?ǜ_���d��9*1a�x�¢��Es���6����	� auoY�:l����tXo�&6�N�sSq넓NЗ�Zܺ�?�%�A�3����m=�a�V�����B���+|a	C�,�������Q�������b����^�:c6���K�2���	E|*:]8(����������?����=��+��Wø&�����՗�ȴ�֥�Fgί`$�.��Β��nAf��JeZ�wm�@���Ej�j��q͗��E���\\�F����CE8"�L�	�U]��z�'�[g����~�Z+��F]��3�!Dؚ:�sl��qD��ӹ�j�l@}o������<��S���v&n�JVnT�̾����0�ZE\�&[�.7�����7{�z�[�W�JQ��Bt�n���$�f�ѣ���r]��[�ҕT�uky�1�pJ�奠���m 2���ݪ���5*]�"��˪S��-����?�t�~��/�����)� ����2:=�3c�����Y����Ml���[ �����LU�_��Q} ت�T�kݡ�{I���(���.��r����Cz��_�����B���K�U�"��!�a��'$V��sਪ�ڮ�◒T��"uy񎫇L�j��-�W� �:����J
�K��>#�A��/x�g���>�]�<]~����z�]8���6i�� F�}�]��`�>R��CX�&�鍪"JH��&��Axj�#�e�H�J�Cc���a�)�ٓ��57�U.�g3Č0ٜ��9��c	�l{�[0���wX�P��L1a�Гe�PNM3����J�$��~86^�0�ݩ�͍q�6��k��V�b��-����H%�WY�+���[���f��M��&����W��'e���*���Ȫ�dֺ�rX$�5��_���N�ZK�;���^�N}`�`5���2U���:U��3\.�;�Ah���Ɠ���t=�N9tp0�J(���jV��3�����f����t��ǆ�啱�v���h�*;Kȸ����Oq�N�~ctF+ ²[�}�WL��$!��O��@�������E�I6�fc��R�=��Z��'UƷ��&1W�hyU�<j���u���+w^)>��Щ�r�	-���JD��o<���V	^N����_Հ�nA|WS��)�hJ�TG�E�9����Ӝ��_��)����lo���J���u��~Wjgǒ�����;�\)b��a�T��zdN���r p��Xw����EOoI�Ճ,.�����2Ļ�TZ��������D
i��������Yh]F�ݡ���1q���
g����F {8���k�ɾ�R�^��6S�2Х��9F�a�����J��
�*��)�w��x�n �Iː����V���n�^�^V�7��"��T4�ܲ���7Z���*��D�B}�z�5���������a�����8!�ɂV���~o ������pΛ�4#J	�p��}���wMh�؎�cP*Al�

���Z�����}qQ	��I}n�GX��'Q��� ��Zԍ����\t����8�IY�,KI��p_ŔJuՔmw�]��J,-����ϐ*�=[U�(l�� H�iJ͈���#���g�"��y;k6����@��=\��9��Ŋ���J�6-�#���Z���8�kZ s�L��I��{ڿ�x5����\Yq��B�)�Yu�(y�G�w̩ÿ?�����|���n|�a��c46���#O�T}f�[��� ��aa�`6dA�P�ɰ�[ƴ��OV%��d�S��c�__4V�e���I����9�WœatB������xk.�m�1�I|���A�H�� ��>}��_�ܴ�	��ƪ��ש-�ow}��b��yJQ����U���{W3	���C9��E��*�6"���|t��_�L\�ι��0^8����P|��n��*]L��`̀��߽�#IE�V7��&�Yq.$*4l8�m��E_�i���������.rE���Db�
�Qa��,[ �7)Z��S3���!O�,�,)�Ε��j�7��\�:�mz �������e{�"꥙֧�P��Pו7����6%����ޅ�rc��K6�t��E�9�^�,@�ɴSǻć�h�Ś�萴�_���nE�M'j��@�Y2tp(S��6��d�&����|�7Z�:Wi�G`�³�@hp�HT�� p��Ҙux��|��V0n��TY�����������K�v"�����w�����!hL%�� ����9�u�1 ��zv���M����oh���1Q���)�� ��=8<�q	�Z��S �e]@QK��.����ns��Ơ�l��>�)&�������xo_�Cep�Z�(�&_�a�k��P��2����פ�"47�V�J��pr�Cq
m&,i�!�u�C�y-Jh�wDmҤ�w,\0�/k "�]nhZ��c�`�y�{�!�<��_?w�SI0�.�C�P���L>�O6�ڗ��è���>V�d�z��l���[K\�W-����.*w��|�)Ky�s	}��j��8�N'/�8u������*�O��m��G_�\&�ԓ-�v�Ve�̔��0�^O�"A�-SA����(Lw�F��r;vrۓl��{����4�-U�q&�8d��; ��B�� �����b��ϻ��%�����Щ%p�"mN���C��
sDPY,O]ST󄏵8�\�"ʎh��cͤP�] 
}����[CTL�U�z��o�}_�<�.� �\8j���)�`i��*ǧ�bn�Ń5�	�'����/"\OB*��{Fw����;���pB�kX�A�06��	G�*�����S4m)�Dz߲�-�й��˨��T�T���7������</��K$���m#=|�:&"<��,����}��+�ֿm_����n|��\�Ǭj9�T>��|��{��*�i'2�ߪFY�:ؽ�ee����H�t���kG�ڋ��o�Z�р25q}���@���22��9�;!�>Faj�D���3�g�|(�>�ak���dŕ�m/��s&�^F�.�B��Ա��Z9�A�������J�����V���ڨ��(���9����hA֠����Ӛ/�D���;QpU!��!����}��hq�ͱ!Y�r�:�`�����y�z�l�e/��z�z iz��]�����pM�&�N������VƊ�kt�	�$�t]|��d��N=�k-�imz�Y	�_��*�\��V *�>����\�*oYTP�K���>��lupH5�j ��I�;uo�@��I`�~8��F�	�#�Љ���
9q��|OW>�&a3����*�B��� 	P5Y�l�~�yx�`8��0	fȆLѠgEM�N=�w���
ƎN7�r����8�6}P��`���N�%�N]U��{^�л��y
L��Ws�K����:�d �T��E�<���γ�BM6Y�ʋ_�b�E���E8�d��(޷���A>\�6P��i@)�}���E\t�(��,2kկ�x�e���:�0�������˃��2����Yy<3����cU<�҈	׸B�H����22rl�Z?=��i�$���Eʝ�,��<V�����cj_�l�O�Y`Fz�� �EU�ߏu��.��e�O�j����d9a. ��+V�ħƒ�����y)��M���u�?ǿ0�� �~�_�u����܉H�>��	�$�7gQ�����%Wb�P��]�J���_��(k�H�R)�٩o����98	�MH���^�����]2�`�K�'^�F�-_O��}�1kϢk/ʢ���ۥ����kdo��ή��~�	Z�)��ܹ�eC��1�̖� P��{Q���ԡW^��Y���U&`���m����Dz)u��۠/~-��=�'^�-ZmY���m�I�1�Û"��8'���g�U����#��2цN�~�g���B�O�nbؽ���88�>��ʹA�["�8��u������VO�K���."��/K��~]_H�yOo��X�C��.�+J1|�i~�ƚ��"�m�ZK�ü���f8�4+߶�K����@'!ݙ��f��->���w���M:���S�G��v��ʒSE^7��2ݜ ,3˰D+�/�����
+���)����$�0�bt�^?.���4���Ż�3J�1b�8�t��T��?���e_�L�ɜH-i���S]s�F�ƹu�0��.�@�����ٚ���[w���9F��6C,�Q93�}Lr�[;�]PU*���T:j�p�d��JB%��.*_�K�'��yT@�Zq?��T�����؀#f��7�� $�b�1�#�0����e<�f1A�ۖڂr!��yA�jr�[�w��n��`�~�#޶�ڴ��Z�XJT�/�~T�J|���W�Ws��+�a1F���N�s	zoF�zH���M���I��M�v�G�x/�k���g
\��]VO:^�[��W�t����+��Ҿ`�:,Ć��Q�;��H�
�@�9뛊�*�J���I���\?b������Fbl�ۣ�%�6��X�'����JM�KV�)o����6��a)����N�v��g�)�t�=-�J`�1������M~	]�eh�-X���~炅Z!�#�)�����PȀ���I![����I���Do�K�h�L����6��0��0㾺��J*L@���t3*N`ݓ;�N�����.U��Kԯ�h�ڨ��(S0N�����\�/z:�G'aL/d�n�
��^:$Ze�[�]H獜W��/�}���ܿ�VC`������f���˚������7�cmRE�7K�:���w1IrΛ�\��iCG����]
Iى{4�-P����(�;��f@8<7��H���Òi	��U��]E�����	���?�n�\cU�������ࣩ4�7�-����H��N��hܢ�MD��s8�ֹ�"F>��|*�{lCU��He��͐ro��n���V{X�f0�x����\���aC?�Z�J��.��޸ވ(,7xCg?+M�.S��Fؒ��ha�]���賧]0	���ƃ�xƐa���<��W��epx��,����2X�WV�ng�m�<�a�-Lc��fF�̄ӊ��q8G���*3G	��ʐhev}��a?�T �O���	�QPm����6�b?e^�*V�������I)��n>��H�u@B2e�/�X_]��M�W�jsq*���JBC�R�i�=���f$�ع/��%H�G������x��M�f�W��lqO�������%ϣL�Y��w�Zy&���;�D��}tm��+�s7}�i�}&~^�%�E�W�l/�AO���`6��(o=��GW@/����.�ދ�a�| ��\(#��AC���W�7���LK�ئ.'"��7��V�4h$,��`��)��}�9h�o�ĸN�?�ڈi��|�1HJ���{�)�jt����<��A��:�9-�S��H'u�����H�_�,/���6�����ʲ!�Qӎ���w��̍�AU1�!���i�u(�>�^}I>�%�+��Aqe��|?��&N��H�����H�6�}��~5��'1�BR�S��6#��)�3B	8j�s��ep��K;45\L���k�ѾM'ev7!���^G��<�^9I���@t�?M4T>3� ��s������1)�y@A�����g�1�a0�\C0[�x�"�Q��Ϟ#-j�Lt�n�]αE_>X�0������.���Ӈd}lX3�|����}�)-�N6(g�2c��@��T�S"k΃ �)i ��'���)�1�rL�J�R�(c�d� i�H�v&��dV;�L�yШ&��T�S��0B���Ve˙���ik�3˸V��f�� �����U���ٛ������~�*�+��$�5�uy�L�]���h����/�4jel��Ɂ�И��"��(�~cZ!���c�O�[O^�\roV���>�𙾋�MD�x� ���i�,z�-����3]���+�����)�MU[`7T]�[�D?�gb�F,��'�&Jt���M�`tc���yLG�$*�^�����A_( �)5f����䒬�h%<�N� c��ko_/�;�����nԛG�b7LT*g��b;��t�a�1����$��K���z&�g�ǣ>ag9�Ҷ�p.z<�b�Spc�t�[
���?0-��*�<�%d�c���w��0-�XuAtD/#�Tl8�ӥF�MQމ�����>6���ƛ]����b��Ͻ8<���q>�
 ���='�v��6�J޾���	�Y}�ߡ������Λw�$4�3.!c�w2��L�Y2H�d�<��Y�k����d��E�I�@.A��vxU���%��4	�����~4À��yQ������VyL\t�+��_�w:I&�Sz�� �~����w�&L={N塾��M�j�#�>N)���K����{4�7��Y<q`���m�Gf"y#�c��R��rl<�+�
؈_)ZF�s�PR�"lQ���û�7i�ħ>��6�(1g6���1�StQ�@�nO��9W	n:Զt�y�"htP��%��֬��JYa�}�F��ޟ��v�۩w���ԶF����83}��T2b�g /���4���9��&����M)L޷�/t���������=d�(�INwݍ�V2(p����埪��Ķ�#�c��o����8_lAa�a\��L�@�Ҁ+ }������( ���EJ��U����ͼ��_��P�����?	J8�R��w"����o�r��7�bv����V�ki�)"��>�<3ҏQ��h���D��ū���gI���6_��:��/0����BXV'�}��g�Òe�/)2$U�H�q��}KU���o���-�d����5"�o��-�!�W\���-i$�mXx7�����ůZ{o�kP��T��`��p��A R��#r�V;��ɣ�&��O��R��&.��,��Y�IxF��#������E��.X�gt�m�B��J�'��ͫ=�V�m[
cQ )�����Ә�z��2j���ʔ��~�A~��T�6uD�I�R���aT����a�{E/aA�����[��]�au$x~³�U�@m���h��r�F����",�¿�=�X�%�����t��Y`8x��+�V�$u��Z���,����D��:�(wA�g�b`��*�:�_
iĴ����ԃ,�����c��&O�]r�+ҩ��d�mo4U���[F�;�ɾ`S��;	���m��Ek����˻�����~Sfξj�Y�1�������H.ߗ�]����O�݉w�3G[w.�Ŕ-tWC2p��+�6�hI���Bw5G���`*�5Gݰa�#��'ѫ�A�1n��W��[��c�wq�`Oe��C>�B���u�ì6"�CH����37"E<�`�r����sҎ�V��OwI��<�z�Cfb�[�����ZK���z�bX��g|��H�1�������7�T�����丼���� ����l72n���{�O��M�
� ��r��>��F�{��
=��[GP���`��ٍ�ֹ� r$�U���)Ae�
H��d:��ZU?�8���f�j��l�<�B@x�Gf��r�����1q/����q����̺t�6�c�^}:r�|�&1i��2�1���Ա�6��d����.���A��W�z�Ie��_l��rɯz�܆���B��Õ��S�fu�����]�s���� �tn��޸ݸ�dԼ��q�l;�_O�,�+ �C��a`�X��RW��4��iW���O����T`N�'��:��g�y�?a���,�j��_��P(��������\��jr}��n��\;D����}���ߔ�E����������[2�9�hr��~�U�{���%��z�����=Uy?��.S�Z��ssF��H= JC�u�~kr�9�L4^�w����1�j.��'6����k�5,�/�`G�CHswva�������"��2�m��J��X����YD��D��cY��p��|�o�D_P$y�@7�xO\�q;�?��Q�Gd7�SS���1ku�+Xj/)�[b_h#	�f�'tCA�Bn'mYT0y?m��'��m�G��X�(��-�.�b���� �I<*2׿(�9+i��l��_���*Ien���U���9| &�"�]-���}M�9�΍EQ}i���:���$��~���/e{�gJG"�o'9Ɛ2�;~���g�>�+�QW����ۿ{�G^zv��G
7��s�e��Ԭ�Y*ea܍J�=A� �V�\�Z��!�	�1�� ׳R��bs.�U$�g�J�}�H��գ��\#��!(	�����̺2��t�o�/�M��`:lH����G��#̯�+�{|�T��������@����� �l�O�?"#���86S9n�R����Ht���M����lW��F�҉�@�@e���57��[��.ʞ}��I�ds�w��뺛z�L��*�J���Y\���#U�n���ؔ�_���O�u�7�1�+�F0�e���F7�YK�ē,�5ĝ�hk�7ܑ��w�����&J�kDN5�k��g�f��8;q(_H��c�}w���(+��p��_����OF�s�DG Y��:�H�
�M>��������X�ѝ����ɺ��������3qE�)"�*T�j��R���G���7B��5�o�_9�Y�G喎���"�y̸���} m��+ja�**��1#�5;�>��T�T��1)w]���0��T\+��ك�\�zc�՚����3�ER��J�ya��l���aBYt!���+|C�d���略�G�BV��c����'�I���`��/�7) F��Q�	�J�]�G�5#P��V���L[L�V0�9��B���JSB&�: �a	'�Ś��rSt#M���c��F���Ѯ�*PC7�D�5�֣DϤӏ�IR`٤�Íg�lxD�]%qʹ��b��ߨ�O���rKi�Oь�`�f����ߔ�g���TXY|7O���TGq�~{B�����$D��i��.^j�����O�E�,�iYᆎ�qM���t�5<>XwKB� �L���T�]�Q��,�|�iޙ)�x'�Oɏ�{V�@d �䆻zT��a�H���0t� �]2������|79�ˬ$0Z{����
׭��6�@{�\߶�ONf/�����r09:o�`�wjE6c��qwW�<Ks˿/GJ])Qa�=���H2J����صl��>%�@o�n�6��v�F��x��R�]��������x=~s��a�i\���K�G�y��7�A�O7��.�K9�l��:��H���TjHDE����	qO1ܫ+ó��
6��b눋�Qe�i��t�.�%|�*�L��2G
���,��(��})B+�<��7X�1XUћ�#G0Ժ��r,�2)���O�EA��o���[^��ŝ�O�*�f�"�ג�
*�L��T2v��;�@�@�3�o�)�n�&o@�=�Iz��z�<|k �E���#?Y�L?�0���:C����Y�u��e�ٮ��Ya��xD�b�Xpx�B����}׬@F�а�mvTw��F����o�}� ��@�>I�-'@�v��3T#���it��-詷����h-��*�Ja�0g����-�3Xv�����ղ����$�iOoR�V�a���vhU�y��A�FeT�iC�LA��6�E%�
�j�@H��W~x�#!�c#xH�u���Լ��R�cu{����BX�Փ�D�T�� ǅ�05��W��~�0�6gcN_�Ӓ��	��B�ex)7E,F,.#i�R����˛dD���h�VǐY-c}?�rj갢DToסp���mS�i�n{�?�pDH���Ta��JC2i`s�O��%4���3a:Z�ټ)�5@�bo���	�
�Uv��b�7�4�X����(��.!3�U @?g��A�*k�0A�Z��FǬ^��/:��F�V�C�ea�/�Ƚ
1j��$��d�,�H�4�]-ƢP&l�4pHȔ[��&�{��5Kab�5��T�P�94=�Ʃ�[EV(�k(n�r/j�-�⪸f�O��Ϯ�uh�&�2��}�m�=&�x�����#��eǉ�;p�?֮H��v��T\���2���Tr���pꄜq˩G�TL�7T���H���}b���;=8��JR�������B���M�6�	�C>��9Cn�m�T=���PELJ.�Q�׹-���3gs�S�y�;������Za;1�7�o$��s}7�� ����΂���5����y�w����^>7~wOf`�X"��q�<H5�2�����Bdq5v����גͶoۑ�E��I��e�?C�=��<(H�齬��\��KE`���� mkQ;�!�c��h.�ҭ�1q��x�����t�=ϭ;����������8���=h��Q�Oq����:��Q��<��܃�J��T��ƣ�|L_���I^vP�c�7�0
��[a}9o³����j`Әۜ��KG5���f�tk�lZ!1��f�n2��.���
,���!��5��!4^��h�����wr��[�xλ'���ȏQ�t��#a���ۿ}ls�:7�,PU
(U�q�k9�+k���w�T�=�i�U`�1��#��-_�A�������&�|�,	�b�[%1oc�WX	B���C�~^����:=����kYæ=����3gbi��+��2�&����'�Zr��%�Ƣ{9//2�ݧ�j`��� ���uZYr�15Ol�ܚ�4�K6z�˚jx��A����Y�ʁD�����A\�:'`)2��ߛ"�I� R����v^�>/����eea�u�NT���e;�mi����%�H�ʮ]fa�ps$~W�g�I�E3o��Z��@̻8G��R�t�� �pw/��ԃ@_U[�{�ƶz)�]���E(�J�l�Ό�|Zl��knc!L���y�-����ي;m,
���EC��
h4����~=�:�,k���у���vOy�X������Wt�DJ��$Āá�I^�bɃ_,�4��}��<�gH)�H��d��&1��9�ɝ���_�0��E�^�Z��s�= %�,b�c�asj���vG�DAҒ^O�
�UާX���GY��,�ع}H�J8#.4(;������Y�s�5�z�`G���OF�5:�c���0�A���]^m*+��Ծ����DJ���j�����Zq�M��rXH_3؊z����#,����̄�!缂��j�J��uBX�`����8l�ɋ˳v���+�
���'�.�П�qZ�w0)'T.�8L��#ׄF��8�U�1��5Ǡ2В�D�o�#,�'��ؐ���W
� n9�0�[�}6V�����Pp>�-p��6���t�q&��?��nR�>񁸋c���l=GZ0�^�cw<��Q���z������G�qK�)ĖN',_*�] rR���C8^{�"�`�<�-�u6�0$�hP��j0Ty�7�:twE��鷉�Q�c���`�g�s�����B/�@F�����l��g��9B��m&��~El��NpS)��L-�(,"��W��*v�����8Tn�K��1>�3�w�Ⱥ��.A��ub��V����fw�6�,�t�ߨ� �.�t5*���(��o�5��3��41Ij�!��
��U�d��������c��¦�PL�s	c
�	�7�{�zbJF���� �O�6����V| t�� LA:�}�*.�������$�� �GݎsPg�8
���Sr��/�dR��rm#b���[޽�HY�B�#)�U��!S��؉̧��i]r;�f�
HT$HY��h�%]��tY�G|�r��
��
��u�.��tIo��.���E2(�h�U�m�nj��I������Tl�^&`��{_˼l�aN�m�~�3�/��_�c�7@%0��Xd�N5��U�(������@���\)f%Z<��C�c���l�:d�'�1�}�R�f����Xߢ.�d��ɮ��$tɱj�҃r�tp���3�{-`�i�3b.��oW���a��w+��c��)����O�-�L����U}[i�Uԁd���
-1r����a��]�o7`j>՚���,�������os�'e�����Y�d�}��qj�a�]�6�m=K��灝^�����@�������NX�������q�_�\�g�-��mi��x�Io���C����#�g�/m��m����ԿqC�͵'��?"��Y�'�N�:x��ꕲ�I�At��U��T��|��:o� &��qrSΏ����a1���w�Uoc�>5u*�4ҋ�FPxΊ�'�2S���!�|nd��	n�����:=�/�K	�t�H��8�@Sn�jt?_��9q9,7�~�=1#��m�b|Ty* ��b{ru�j��K�Jk}�����{u���a�Xcxc��v�b���ؾػ�����4�O�+�z3{�APW�!�0��B��!~�,�q�X��j �~Z|��Ó��u��ĽL��+���\�^l7�=t{��hleXq���D]O�Īx��?��_e@U/=;-P����r���1BO;/�Z�c����oa��U������$�'�MD�2(B8�𩰕���9 "/��I�kA�ϟ���㖀S&��k3ou`�>�ǯ'*��J�3Po������2�c���k�Ϗ�Q���̂�咔Q�r�z���*O�}z��9s���l�C ��R,�L��r�����Q��.6����H%�֘�֟�k�;L��u&�xpت��s��0f6C�Y���y*���|C��3I��XI�m7<h	�ϟ�U���C�ܙ�i֋"ƻoBab~d�Ui��h���1��eP97��rk2��J��<��On_e�SD�V�c�ѹ�t�O���?57QA�Ň�R��8Y�o��)���R�|q�r��V��&Q~UɉH��0j�:l|� <)�t!����G[TXa�hh"��9������,R G ����9�sxY�ˡsb}��0t��8'�(��\6�Z��R�Y�B�a#�
<6��y����o��_�7�T�|�M��bg������!�K��wk%�>��t�Eq��*��K#���Px�_T��-�b���}�]�VϷ��olo�U������J��Փ�M*��u[���<]�S0�F�Wp��r�w@�=���-}��mEcc�BȈ�;��HGd��@#��I+�В�h9-��?k�ԜryQHK��^�0�:W��|h]��ty&�ar�u�Έ**iɽH`�/u��oĘѓ��a z�qz��e�6�NW(�uHp]}�6ʫ�y��W�nb�c�a)i��Ow����T)[X�#A+[D�J��;>
�$r)�OH��"�%�c9q����`m
S�aU�|�d�_���,�b����O�!B{ͮi��R�yF>�8�oW�}��AJL�f!
������+���ޯ���t�Z���!&�wy/�ș �ѷ�����Gv\
 �3���(�e|m�S���7Sڠ�}�-)_�9^��h�Q���x�j�-?dd�������G�f�t�%�v�;ESA��:�譒B(l���[+�q�.�m0��_(:l����cUf�6A!�7*�s��W���c̕Eän��$��dbٱ2>R��qݛo�5ٖ�u�z��'0����K'X53�ZZ�� ���at/
���F��"�JR4l0�*:����<u;�αL8p$@ΣRh�Z� ��*K-���#���(tƢh�v������Z�D"e��6������h���"�}�������=7�����H
�_W︫ȹ����BG��Rr^���I]F#i�Ր�~���-H�xu�?����R�J�� $�=�|�e�
�I�
%�:�[,�c��Ė�ϬV�ׂ)�ᕀ��G�ۏ��6�qc��!��~xo�#�R���+��K �����i"r���gDEC�����6	�#�����3Tfo��)�s1�yI�K��*E2IEQЧNi)4aa?9��{�a��������ޣʳ��u1��D����b��n�CSs��$�R�;�I�P=��ސ]�m��t|��hnM��ί���n�e�M+H��^���Ҍ��n���2��t�{ד/a�C���a�=��e�Z~7��s@(#��f��I�Q����v$��m�I3Y�A��pq���W&I*�s��Bِeܫ��ɯ�Ê�ik)�YU�����+��/!�g�=� �x��0���g�B�zΣk�#�&�:���:�Ä���9��LP��&>�w1����g��-_���Pb��n�V �����|p�V��I���H���qQ�bNI�$Ω��o�T+%җ��5���!+N5<�nY
��RFD2{�N`�IimKP-�-� pS��ȽRfݐ~�`���J��z��dPx4`��g��U-ʡ�����I5;���9 Q0���������n䱂�$ܬ�S��%�c�}dXs����he�-�,O�a-_Ӧ(�����3@�:Zus^�H�E��$k�-Oа�h��;JxU����-Җ�o�H
5�o�m�����@�b���=����y��9}�Zs���*"�N�o�Y����Nx�Y�1��Nz.�׎wz�^�!ec�}��R� ~j�u�M���0$h �uv���(���tO����V�1�9��G<V.�k���G��?T���o�#s�edq7�q�?�IU��D�5ޱ���I���#��V�e��Ǹ�;�`3_�S�G"s��԰�B�)��G�@ǝfg3�ξ�����'�g' ���8^Y6�Yc�d�;�)�PC�R�u��x��;��h[s����ˎ�|z_؇��h�cl��ǈeSe�8�,����|[lF��?f�S=��Tn�4n��v����Vu�eA�<^����z9���F��#t��[a���ߚ�ǎ]?lK:������2��1YR�&�Q�+���7*�º �	\�����bӽ�
��ࣽ��eѻ�}a����>u���7*C���wG�����y\+ٞ���;�3���ᤒ��x/#�)Hխ'���ZJ��mL�aY���$�	Ϧ�VH[|�����n4n�����RS;Z�����}T���K!:�
ݞ�D�����"CB6���|�1���@������ �͡Tb���i/���
i���|I��±�|E�K���� x�oag�m
m�m��V�j�G<S$u=03�]8���y�p��qc�=.��"��x�R�MG��e��ZHMA�kb��Ι�s�{vH+WI�?EoU,g���wÎ��m�1�Q��уu>�<�ˋ�0s}���kAJ�ݽV~��)��ʥFDȆx��F;��$���wM����U��u��Ǧ7�ΨD�w��>�?���rl.�=6�⼅k�o֣+ Qj��� �f��-�拗��u)�_���ɃKE�#���Æ�}�1��6�}l�����y����i�<W8o�(��X_n3:�]c�\�(��R"�,Luő��n�[+:q�~�#!3Lt~�w8�D�����p�v)�}~c%�x�C�A|⥑���*B���J�P�W7��,l9�x�%��z�ǖ���q�}q�`��D�y�j�[O����h�8���zٝ�AD����P�6�I+�1��9�@���C{��92�b>���>6�x>8���%�Վ�Cy�'�En�-���cA�<�skV�@�Ae">���*���aT<)>�V��4t
�u�HFe p��d����/�̆�@Y_I�x�6��{������RO��hȜ=7k�bFQ�L�?w4̈́UH��OO��Y��?(M9	D�;���]����{ ���s@\� m����	�6�AY��6Z�>h�d���ʲ��*�5� �����u��{?��"D3s�Vxa�H��̑`c���RGEy���r�e��'Y����l/�*M�O��Kn)xLo���q�jE��IKl�>`���t����Jm��Cw�l�v���ƒ9#��8��+��I1�;k����u��%e/��y�S��b<�8M:g$E>�[���@3�urp�e��OH�ݷ�w����=y�������ޝx[)�c���b�D"�g-�Q��� 7К�sE��0���*�Z� �N��x8��ؘ�A�:�SZZ���c󵕕�{~�K�>lCے�p���߽�N%�T\���v��w2�1Sm-j1�:1x2�JZi�<3���:ú��õ�w2�\ �j�2�G����"f��f�+Dޢ��(���F"��;h&�:.Øw��$܄V6�Q�eߝ����K�2��G���	kF��S�# ������Y9���!�{{E���U}�¿�.e��VyC9S����x|WD�AE��\��Yl2]:�V!�O��{���u�50��,��,(_��=�!��ϗ�1uof�[�2�z�:�*;��$BFr�#Ĳh�"���gcF��ή��J�f0�:����R�5ȵ�Z�E	j��?nXaw�9��<�=���e�#Fi_l���}w-�"Ȅ��ޭգ}���E��!,޵�i��U�b����Q��q�#xMg��1�'�\�*����,�}|o�_�AoT�� A8����K�aC�&ꐨ��cqR�$)�|XSy3�g��
��Lٟj�Z]���غ>95+u������s���.]D��P����6Jj�q�3��z�	+���XQ7�e��Ԗ}�D���t��K�MH1o��X9�O.�ƪL������dXF�.H_}�Wʳ�:$V���:�=p-�	;I �|Y�����ܕ��\�.~Zϓ}�6�2_�u�����a���?�-ó9}��M�Rr�J5�*jMR\o�������L��b��ޞ4�\�E��Bԭ�\�|&^�-1�'���l����˂6���v��!���4m�c/]B����E� b��f�����b�L/�='�NI��0���e1�$��t�$E�g; ;�[��f0r�mb����A:�>q�L��^���R�䏧�\>	-��G^�� @�W╍�3���X���\z���[�%�Ɋ�&gÒ��ƣ��U�@�o`�A��w��5Ҍ��[�`5�R]�f`�Z�x���3��@(>i���C��cG�1��] o�5�%�_� �p�dM� ���Ɉ\��z
��(��/e²K��1��s�e��p��dh�DL�N*͕/:��ʈ�b��րd���qQ�`P�P.�f-r�b �Z��9�B��pj�	=��5MR�����(���EW��^f�E��ȆwC�"}������7bӐ���+�}ř�5B�F��r�|�8�={�;��(l�D3r}w<��.K,�^U	e�5y�F�h@S�)��-B��1NůA�@΅��t)�[#34F�SK�^4D;�"�+��a���}v6&�0$ �:��P�A\����k�
(Ɂ��u����ri�-�~�,�ǈ&�Q��IK6�ZnM�?ۥ����X��C���B�\��7��3��v��b�~?)4�r��6R�ȋ�`֯Ǵ����mB*8s���F�5�HhOȈ�]�1%0;�L�w�su|�)���}>��m��l_o~Y�mF1,c|�.�$��Bb��j/�%-�:F���lW�ibo��eW�W�*[��I��;���Sjx6�Uݘ�.W�+H՞�՜��Pf;^;�b�g^����4	5b<�dLg��5�rz���`g����z�)`P?�L>�M����"�K�[Q���l������x��.�uK&�?#�O�R�4p���U ݋g^7h/��@h� K,�o��M���t�F�����
�.��ѣEI���	3�	�_�8挡��|_��� ';D^�s_�Z<�~7��+�*���'��-A����E�V�:>��(�0��Ϝ��Ѣ�4�p���`C`I��5(�g	�1i���D�Հ��a5�K�͂>��6�M`��(b`�=J��P;g>��k��bE��P�f���:�T<�e�)y�}�b����@/�z�b+�ǒZ9oo�V|g^���1M џ�Տ�־L0?ܥ�H9Ѥ��|���������\Ъ,>�]6i̔ɍI�i�;�Q(���>,�s��̿�$�����c�O�Y�KG:� �Ӗ՞�%R���l\jZ�@���Ź䅁�"��̦�����O�X�x�>X��
D��Aw����P_�&��3���8��&a���Ѥ�!��/��m�c�[�q�{tIL �N���[�]``��M`���[n]�A䗟+�z=	�v!\S�g�U�΍�%+e�����D�^y�b�b�{hhK��)�����E�'k4�Z���{�����=%�ig)���˒��I�*�@��t��%��q����o:��tE�PK8GÍ�v	gU
��+��5������㛱%b`L��*>v[�$o<G�=o�-�|4I��Y PXdY����V�N�F4a��5�D�M���+�®|�ռ����do�tȒ$_����`p� 
������˦�vN�jȮ�JF�͢Oϣ��PRrp5iԀߝ�ϣ
,\�: �r����A3�I�1�/d�q�8}1��W�n��|�1�5?�;{�g��;�t�X�¤i_�`�@��i�u�D�������T���ͯzfҿG6�R���{{Y�jNQ�BeyCWr�����,�v�f�W����-W�.����e����W�>�=����������Q�R���?��!SCn��O������4X��8��S�Y��oypC��?�,l��0�b�4�wB�lM���x��%�L�]Z�_+v[?��W457S����	�]�7k�����[1���#�q&4N��`�O�T�F�v��KB����&i�M'�}�9Yn!�^�U����'sHAo,�7�
��]��ٶHjۘj��|�N�(~Um�����s��x��f�JbU;mp'�L��������!~���=168%E��q�6���[srd�.�b�Aʌ��D�O
�̦1?zPh��o7�V�ݥ��ٽ"�����`��<���c�l�`ʡ���DȺ��<b�o�!WI뵹`��gH�\\�n��s��d�mk�G\p�q�ŊX4WX�q�5,h�s�萗� (��z�OÅ�ABXw������Xr��m���!���.jlD�qTt�^�nT��ֹ�!��HT��8��vQ�
�P|���ϣh����=B�.�������ǾIy�#
����X �;o�%R� �����_�7�|=��N�A2vw��W�m/5�q{�(�z�Xu��ƫ6�?�~�$�t?�F�8��7��θi����`d�:��Z�}ɭ�m���?/��Q��D��缱�����a�@Io��x��65��Q�&�zYlmG��:�5H��=7���zƺ�*���>{"=C;)^���B��y�D@JtJ���Km�}�e���Yf�e�N`)��D��֘����a�,��e$���}�G+��z��S4����zu���1$\cn~�#�|�1=E�Ƙ�Y����叏Y���4�f�I0���u؍64�}��hy�:/��t�e�I����5�$�q)d��P<�Z����pdn�GP��9���5�z&?����AY[��I�g�CL�J�\l��l�֧�����?o$��h`�2�o�Q;��.�X;��nN�fwlSnZzIw���d�yk��Y��O���p�!�@�$�[��\�	{�i�ì�ȑ�R@��ǻA��ip�a�����k��";\c;�:�����0��lX��䄦U�	~O�T������r�x?p�2��b�=�����h*��Gc���7�܁}���4�[�=? �C�Tj���t���7/2w{�@N^_)�wsV��72?)��L�.�I�G�d$^#���5D�C�,V]Ǟ�:Eit�b�,���3����B�Q`��0J>xJ�XS�Jl��"j��M<�JH�Ͼ���Z�@T	\�XtV��U&v�3�*��k}gϩ�h��������G
�/����~E�Zыz-�nȵ')�4C�~%��~�\�^·���Bp�"�I3��Js�WC�?C�.L����������G\m�S��+�_I�xw�$�ʵ�*�F������_K�I�g6��ņ5"�FJ`����`�6��6�ĩhɭgW�y��#�=vdA�E�\��8P	M� �� �5p;̀��;��1��@у�g�tQ���4Ivi9� ��GNڎiv���I;o<-?�,��	' EK�|P��V\{l�1�r�-,����:���N�C���b�	e�|jӀ��&�����,� �g������� � �B{7�J�*5��Pd�W&g2�3d���l�Ѳ���C�?�i^��3S���G��[�"��D�MŹ�D�Q��C�Ȉ�K����q���3a���C�ʦ��F����V��[iޜ�9��C����0<\Y��S����L8���*,t.�흡�y��� ;ۭ>k7��*�A��5�Y�<�Y��Q0�vi���8ϣ�M�����̪��A��x�	��T)�(�\t. 4������cn6^�b��ֻ�f���yi�@��	�x�P ��/�2W���m��o�\y`�o�Ō7W��5:�m�<0�ҌII6�jfc2��=�h�k�R9sˋ�:T�J@��~L�4�erc�#�>O|u����A�n�Y�4��"T������a8��͡�׭T�:E$�{J���䦊yʫt�*33��C����#�55����<a�+K�_?�����c%�O��x�P��	̋����했�#��p�EhN�G,X�R��Fy�CN��Uvg#ۑ�����#K�A��:��))ceD���L"f<GG޼@ʳa�O	><*
�kK뼹�hR �,eN�-EV�����c����p������z�]�A��jG'�E�DJ'�
Ze��ܖ��[����w���/���~��JzV��;7��>�N[��.��fa�5����A3p#�~vsY5�"\�P8��]㩬űRAj1�n
2��/��V���v��u���Zn��;�+��p�_��@��|��J�(�*q��rz?�&ĩ��9%�9�̄��ɥ<���w�15^ �̍4�'S0�6�&e�KD��*D��`C8ӯF�^QL�@��`܇�T��Vy>�z��L�.�lR���=�/��gi���8������`��p��s� ���)�0��)�|O�uu"���A���tҦ�fChl {�e�P��0QT�l-�<7 �@���M��6�T�K�]^�㌳@�8tiP�_ŘE�R3� ~�mDb���ӵX���˪���n�Qꆹ�p�ܞx�s#d_�Zfg�S��
pe�k�@U]�]�܌���?�n6��P���k����3���1fO��vg�0�=_i�Y>��tq���>�9�U�K�9��ܡ�c�OZL�ƫ��ڄR��EW����c�gmH���Du�dG�K
6]e�V�x���1�9���玲� �ȡ�Ԃޚ�9�/�UWv�7N�қ8<|�����cV'(�_)�DF�R�i�%-%�W��"m�[9�=1�������h���;6�Gm6����V3��o�	C�VUQ� P���b���f������.���mۙ�2G��¯�g��A�]5W{G�� ^y2�**3�r@ �H"#�@�R�
_޵S%s�,C���ߢ�[01j<D{u���Ў��#Mrqq�m�d��8���;���[��{\^|J��jW�+��������ޭ�Z�؈1���jq���η�[aqF���(�KV�L���(IϢ�m����)X�d����uN��Ac�'��+Sw~���쬾\!IM�H�Ϩ�b�J\]ꟍ�}��M�d 4	��W�K�.I]��(��7-UZ�\���L�jvs��.����|���o�%a�/�C<��W�}M��-�>�&����x d}��3��]�o��ӭq�҂���$��
��nx��P)�#�睌v�2�D��@i���+�<)M����ڍ.Xs�Q'P�w���V���?��$[3���m�����_�ܓtJ�?79�c{��(q�-Ќ�^�ja����B��)
pr{8���%�)�z18|[9"��5F���4����n%N���܏cQ�=��hܲ{�@�^q�U�Ӟ,)Q��5�TlPE+ K�'���Ѡ*�&�Z)��n�E��t9��.��C�u�X��L>��b��U7@����� �5��.���F}���!��)�����OL\Y#>��K�A��F0��I�R`F���yd9�N��WD�c@T �}�I������y�1,�2C���ܸKmV� ��pvGz(�巧"0/�B[(��+.��{�_G�R�Uh��g�J@���(��AnGP�B�q���]���`t/� �N�Ǯ�1T��D2[ڳ^��|XX����]zQ;���ۚ��\ �5�(�����hP�mAj̪STI�DSE=C��S2Zě*{�qe������5	��i�"�2o�qSH�El�t����3f��`���I�bӹb 
�H�{L�Q� }�}�U��ņZ��.���?�{��Zq�eO�F���Y��{�Rc-<�N���������ܹ6 zF[IZ�8��l����>{��U�R�"���>�3a���4� �&|��e����i��q��F�U�:Z��B*+�4CB矄�|J�o�)����Hx~O����f��KSO��*��j6?/���\���Y�P�Q��Tw���j�a7.G��f�?��}�y;�퇃��82��r��D��j~�_G�h����m��~-����`P�X��)�o���]t�,��Y�M�U3�Zf��U���t����eM����k͗��<%|Pa 3�aO��
	�;��O�i�c�|��bg�[�_7U'����W��x���C��'�#�.\���@�nd�"e�n�D���
�����Y��o�o��o�>�C��5%I���0�/ @*�:�M��G�,���~�ޭ��}��\N����\_���1�܏)��07ƃ
�s����]�د��rF\���p������:���t+H�6b��cb��wH�a}c���\*r4��%PL�-��6����#�^�� 'tqʓ��ռ;�>G���%<v8�7;���|�K��᳣Xx����G��F�7��<�c?/���'�}w�P��a�4݁��7�ܕLv��D��mc�p"��RY.�K��Jb�ws���z�&4�yq�ty�A�&>�"|x���;��|���W~+~$Sk �'bT��R�ĩp���=�r'��Od A����1���Ǩm5�"�l�f��1Ԛ��]�'�'���t�*�/@�� s>Ͼ,��N��"@1#��N̖�9����ݮ�΅\��+pDs�I��p.4CR3���X�Q�B[��m1'�A��>��i�goc�
{HrD1Gb_p��!�<ĕ+	��ɊY�U+�֮�.'I�}hD{|ː���U* ̷)	��ͅߪ̽_���4.t)y�`	L1qN�1�����=����o�z����_$ӭ��ǝ��`��s��($�TYy���,�ߗ�����J���T�WU�u�`2M��EU�e!M!`n	t��p����a�j�U�oB���Ƽ�b���Y1���^Y��D�,��,�5������EL�<ci�e���R�,�?KW���X&UH��]��%Dٖ�H��u�1�(/����,�0%��9^E��-e��nO���l{6s����_�"8�ո+�N�0�#��3����@��\b'Z���s%t:�&X�|�^p�_�8�=T���Rw@�$O7I
�2AZLLc�q��!�IE�b�nw3��7ێ��L[��2�N	TT�(����5�u��i`=J�5���m��n�^�A��a@Y��{�42X1��,������I7��-;ټ����X(�{͒#4J(��h���dN���I̫*U�{6�MHH�_R1h=�(͂G���\��T*V�?�l�a�ax�q�c�¯�Z���ʷL�E�6�Je�l㖇AS9K�H(W���C�>-�ة�J����AQ����!�e$(^3�a��D���QG�9,�U�3#�Mk�xZb�g~��1�fSp�d�^��{�A�F"B"�p��X��N*����������m̩B�s$b{���}����d���~�_D(�J뱏.��4�@�M��D'yPc���f��e2c�T�)�:U32�ւ�����;�Kgs]SnWA�i�8�������.3��;Z��a4,��Z}�fHI_��b��\��|�=���0�rp�#qlS9����&O6T:W,v�Ղ���yg��z�H�3���~y7�Z|\��Pu렱����D5��/��)"��N*�n�-�&R(�����,nt�G���R�f����q+��򼨴Ԁ=���ho@�U&�u�s?d)����ƭ+5����k0��"�����w��F
���7�ҵS�
_\9j�ؠkv0���b:������K�<2�=ۍ\fA�##�;�a*�*��[�,8��ku���Ɩg��8s��C�Й��A����@�����-�"�������>���f9:D��Nqp�Z��FZ�E/��eTR7bT��{.F��-dЌ����m M���/� ܡ_!w���_�*�LQۑ���Q.� wM���0w��_.Sѱ
�̧�N"`��������O�,ٴ���QbE��P�5�!�Íw��X�M@]h/�o���C~Fy����:cXnJ�=7Om�G���iG��k�����(W��h��?��2���㌀]�=�wD��������f-W�9C�	#}N��pn{�m�Z�<��b{oFy��k%
ΒC4�~�}p��%���oH0N$>��͖}=+�1�
/���v��
 w{!�C������L�A��+��G���ȇ!ޘϕ *�u�iU;H]�=��.+j�ޙ�9^�FDo+r!k���Q��)�N�R�~E:�SI_�x��=���JT����x�>��$BS�wq/����Ci"��?3z�ݪ��R�vg����r,��m�#;���{ZEO�%��� G��l��ͿT���d�j��=;�x�x��	b.)E�̺9Yٱf���\R���2Iq�L��9�P��w���t���Ϣs�6�a*Up��eT<�Ժ��o���M������@��	�K�vB4��r����}b�ّ��/]ݤ|#��1����&���vD�a��!Q��!���������zՅ���Fs�Q/Ee�{�C0qd�.s|ٱ
�����h�!Xx��`~�d)�P:X\_�|г�d���Ξ�,�f� �qe^�����U�j�l\�VV.(*��d�y���{��b�.�^�.�\�Yt����l�U��TJI$&�9l�K
�3k���Z|4���'��Q�N�<:e�:!	v�3 z��a��t��f#_���L
F:�D a�� ���R����@Ì�#��a��O�26�ܐ���u3"��?{ �.o�g>l:m�k��6�ۿ�|�_6zW�'�y��V�� >V�����N]d��!����q?,@�T߀@f0ݏ���i���!Y��EC
X G1h	�
7�O�o�FK4���fhٳ�$T%��S��4���?�3q�����q&[U�P�@�֢�L�ʯKDАI���By����Z�Fc jE��#�J�ۏ��q	w`>}7U'cvU�|8x�:]z�K�1A��#n�<E�u�3Em�J���Z	h-ހɎ��.rl22���Z����CI���M������N�/�1�52�l���X��_��G�I(�\��Y�d�{�S.�*�̻0)�1��]�C�{��v�
����Q�����s�!�T���h��A�dg 3u��|1�� �j�u��z���{�J�A�]5 �c�JL���9(���T� ߙ��x�h�d�����5�:�J��ՓmwCC4��I"֮�y��"�K귾M�ը��8�F�j�#����f�U��Z^���ކ@M7�+{/��\�\%1�.|��źuU��T���O�vEӳȐ�������>��0�S��9`��VL�/��mYb��/�2F?&�዇t��P�Y���SAd�;���l	�������,��|����t,m-XR�p{i�+o��s�s�S\)��Ϫe����O�}��)��1�^E-$a�4V�陘6�Q�4|���{�{xY�4a�I��~<]���[�m/��Xu���$��c���j�ZB\�se��{y��w�8�􃔅xWP���z��4�^5k��-���N}�3���EW��@ ɑmO���Xz� ��Mml�.wX1��A}�C��C7�'��ln���9�Ň�(� Kt�-������q���T�m�&Q'$�^a�`�>�L��XL?���+���r�����B�	�V����d�l)��+̜�}S:�u��c#��8jޞ��.p��m�9�b�	�] n�!9�[m���%	
85U
V%[����W~|V�,�˾�T�4�iq+Y��~ť��(���[����)��>f�P�ut{�T��`�c���Ќ;�ݽ��2����?��E����ݣ'�!D�D�oۀ��2=� 
�`\��B$T�]�;��|IE=9 W�{���ͷͥ;,��H�])���K����]	ѐX��d��� �)9��j/�D�bW8��2����p��S?w�1�3v݃z�D1�}������6x��� �>툐1_띝�>��^���<:��p�R�!<V8o���q� �4A�xy��goEix浦.����H��m�i�1jH�c�=�◙z&{\+�~�h���8���=v��Α�ZN%�@(h�s�~ �����8d���kD	r6&$��e�\�4`p����饚ɘW}���	�:�]��q�2��-�ސT�&g�?>�>����g�	jX��H��[���É���Y~��&Y
Jʫ�4�P#;ӣ��Id(xBrH�ŀ���L0o+����#�~�>�er��2�R
�)�z��V?R��g7yZ��o�-�f�]A1W�z������%�T���K�3�m����;�Ā�0��2P��R��so4[J��G�^bo�Z�}��[���	����8��op�O[���#��w*$�1�3�u�.�^ �'��:�̻��u��t��!�Co�-,Rw�܈ه斨EnG�I�7KqjY�b�Rb�ZI�������Ҫ�
���c��!�9�>(�
��T���=N�4�(��Gy���f�҂�YB���鏼|)������Z�?�%0�^܇�%\�� ��a� B~SI� !i>`�]ޣ	]H�6,����#�s�l@慹DU4�IFŻ�_�8+`4��7"��ȧ�CkG��㽷w����$,�_���ԯy.)���\��L�����mTqƜ��i�%��W)6�\2��^re�Z�(�Rp��E%U�7�f�N_���/�c�/���H�ј��T���,*e	�����i�Ȝ��=�M�:Y8���I��[2�)&Z��̍�烟�0��^�9R~��fw��W�a;rj�xIQK`�)::`��v�'�PPٞ�� �mGF�_?j���]%=��_YZbg�|ȡ��0���'KU�|u)�cm��T������]l�Y3�G�� b@��[f߷�gUR)���h�G�����i_�mR4#��O0 {0h!��o:�D��'9���	��F$��� _ ��Q7�|΋y��A�ե���Po>D��٩�|#��<��ڵ�v���#<Y)=9M�|_$ʊ�X��H�>(Y�N�`q%�n��{%�>N�zEm�����p`�����>�V9�V	���ѷs>��p�ӓ�~�<����M܉+����V,���d��q!������rj?�W�����ާ
����������y=n��?P������P9zI���������ŭ���l{v��:�>Lc���К�XLĈ3�r/��d}�5���a���/��:��.�E?H��<�[!/���+q_6��@}��OBμ�}s�欁5��D���Q�q9I�lw�e���ҥ���u1�)ߛڵ�v��G$��m�i��h5_$FضĢ�8ؑ�"گ�/t��Q����È���4h7�>cw����E�(QXA����r�#�W:��A��'��^�����Y>|��hV�L$bX�Q8��Q�7!�ig�]gr
=��0\2���$��qz:��@���i��h���U����/_���y�0����Ū��vTR�Y��\#GD@,��(����n!^���~�����*���ݾbW�+��)�YW�5����i��O�g\)���I��F���@�Y¤���"��X�Sk�+�8&�EJL�?b��Z��P�>w˚/�8�(t�'��h���ac,N�?$e�T0"ɀ��ό��[����2�N�*��X};ɰTA�\i.�s@&%�갋�
Aw)낊�yo��p�F��`a�)�s�����!��͊t�BK��5��+�.a9��@�����آ�w4���=����{�/��e��(:���+��$e8�1������	�P$��Sa�ɍ��3�f����X����K;�D%����8%�X[�,¾�3� 4��3��=��qUB���ɰ�;J��Œ�r6 �iȜ�鵬Cy J�������yy!��Cԉ���E-�J�i{3K� Q�+�L�Vz��-�G���&G�}E�&����/��O=�9�#NEY����6}䇭��\��.�MR��O� ��WL\�H��l�X��JY���P�#��ǝ�,�L�LO�5�Pp�;D�1���8��kY丹G#���,n��H_�n'��W��\_F(&&/#[��T����㒮�l<��_fj��,�t�� '��J��|MC����Ҫ��6H���t�Yk�41�?9���q@\��[ՔY#is�`rہH�f���Z�ihM5��\}M�UC�ٌ5���^������f�m:$�m6��t�s,=%�e�U1ĺ�����\��t�'��^�j_C�|p�'�+�~��S�n��l3��A�Dl�Sq&�{��Z7�M�MZ.X�$ӄ��{O8��r���r�����޻��n��r�Th8!����QT�fNb��#��$��6ϵ@j 㧌����Wk'Ǧ�G�}u?� '���zk�|6C�r0}�e�t�� �7W���U�	�ь�r�I:z>Y3��P������KL� ��oWʵvu஍�l��H������C���%���a�)��*�N�5��`]��hT�E��`�D�(�����h �~�[�oҒ{�$�iZ��0��2�Օ���Rl�Q��ip��-�5H�m�l���Wu-\t�ծO} ��݄�D��`���"��u��^�؈�3~�M&bV���f�L��bO��&�')�ì���[�$\�O5�\3���&�#���L�GbE�5�=KL�$qP��z3"G �X�,��')�f*�lZ�M��-{����Ɠ����;2�f98!<°E����~׆uZ�K�����t������MK�b���+�����%e�;��O�0�����V�`��������H�)�G�v�U�;����DY�z���6�J�s����|_�g����.B(�����!�_��7M���luW`*tI	�I�^�����{�~e�w.�C�� s �e��g'�S��g�/�7�R��1�m�\�'��c���<*�'���b
�U`H[�
*С��E���>��,}$����yR�m�!�
X�V�C(�ּ�0�馷M8�M��{$v@Aϔd������\-�4��P�|A��0�,�ԅi������93G�X��e����<ʭ��פ�:V�hT��l�ͨb�ɮnT�ޟ`�J~S����v.��1�|���w�.�/���~��и�&��'&�3�xQ��P��z�]'���A*�T���C�>���L�,���f{�V��NU�Us?��eN�M���e�_@6�gVN�2c<��M<�r��{-L�5�C�C=���K�j���O�l,(~2]پ���U�3#\@'t4)d�ܩ�������`��o'I[ҷ��s�U�>6�LsHZ�)��^�z��m=.����nw@����H��f���zD��}�{T��E_d<�D�cT��P��bw�8�'��b�#$	<	,���Pn�u�4�MD�sP�b�B֪_giz���ˍ(�޴��~<�P�'b�oL�``�T{S�K9�:��j9�Z���k5�@8Y��!���?���@k���`�h�ld��{� �W�n���������FyPћ�u2��&�LU��nQ2� ���� ��W��ձ����=���&�%P�����T~������C�g��b��b�e��e�� �f�����kfJ�f�˶��=�
8A-�C'�r�V�mλ�MR�A6�"0M��7�H��)חuT�-����BC/��T�"B.f�
H��{�o&=�(�`p�O�6|!ʆȈ�+a��@i��X,V��0d��`�M�,�]d�+��px�v���S�@ڕ=��H�o�(��?v�j��V\�:��"��M苬E�B^ނ����=di*�i�͟�H�U1ec�ލ幝��{��dJ �M�Z�h�qR"0��O"�[�x��K��,{�?3�FH�:~�� ��k-s�H��=��*�� z�W��Zgw����h�U��sX�����G��{��Dy�&l�R���^Nz�Р���ג�E���)�Q��ۄ��M����S��9��f��s�E+��幆L���S�Y�S�.�����@���]C���eh��2o��������u�7����������0��js�;�URt�ШU�e������H2!��~�����R���Xdb�5�^eq�H �>��85�;�r��٤��3|�>�M,G���iJ�D8���J�vޛX%%��?��<�t|�$]�Nv����b9=��<ūC?	��K�j-�+�ץ[ $o_df�k�~����Ge���C�lQ�}�gR]a �:�_���vv$){��u�0o߰l]�=�4�P�����-��C���M�i����c���O\1����v^'o����O
�. ����@�a�KZ���[]{i Gd̊�&���A���z)��U���cXo;z]zQ;���a��f�A��љ����°��t��nF�"�W�%V����.��_^�J�d�g�k&y]��������t��e��\W0�bb��>R�ۛt�@�Z�iN�_�(�"Pћ9�?��Fk��q�ͤh�ƍ��(�#p�X'6����n�fDO�ޤ�ÐS`�<B?��t6����Hx��oE�"]�MsJm��U$D�~o����1!ј��%��Qc~�E���p2\0*/�a�h�d �(g������D�B�#�r�z>�	����!f��y\q�O�"�#=�)�od�Hꍩ+�S����+Y%��G��Di^�+PYY�v���{���R��ɽk�k��G׬�MnqJX��nP �0��9��l�ǩU�-�(D�o)�N�U���g��/E����> ���wJ�M
J��G�����;$��q�h�s-�K�ƍ#L���r�n}ZUv��Y$#�,��6�ʜ������P�Oj�pT�5{���5�*Ω����V8p�5��a:�/wB�o.����"o�%�RlIC�LGݸ	|#�v�xil{$��c|<������}}2��I]!XW�A�:�����8'�n3�lau�
O�m&[�O�T��?�ǫ�c4�
��������_u��O��q�N��B�"�x�C�}���
3+�G-a�ݗ��`�i�~s�8�����¢���b���mC�������F�U��?��A�����ba7O)�)����"#�9��V)3�R�ݥ�*0�6��s�q��3R�w����H 9ҭDJ��L8V��,�nn%m�����t�@$tw��7�Q����/��`���|�h��&�@u���KW����$Sk�7��j���c��կ�����:m�ήږ�~�������ЗsmtF<�@���?��V�d���C��[��ºeԗt��g���;�o����7-�\�"f���}V���@�r�A2L^X��)A`v�E�8�$�ԕa�K��uc{/Y����e� ��$.Iu	��%��Ԋ��������F��� d{�.�?�8��UR8����ǹ�`��ⷿ�ڈam>����'�=�/�H�{P��&�o��C�͇�� ,֞v�i ���qm�����``a��ʜ�-e(�!������V�7{=Q{�Bj���P܀����w4�9���4��~�O9��#$7�MT# �"
Yf�K���E�<w~r�����I4�i�f(}|XZ����$��n4즽�̀���_�`�I����6>���ڊ"�g�6�Ԕ�� ���l�rW��v:�{�ݜ��`�H�Љ<�^
��
��Ed�uE8?�; �]��W"C�����p��>�d��z]D�`��;0F���>wؠw�#�Q����{��@��b*����]3s�؏ D�?%���Bٯ���!j�w{���{�AE�Q��|u�p�N��<� ܛ�΂�u�~
��U��� ���ˉ�0��T�F2���o%�M�`<�&��a�)�̂7����-�c� Oc=M(�`9�Lg�q~�B��ڹ]I􏵐U��w���=�㠢��>;���0XyY.8�����E]\�4��9�i��gr����O�#�9SB#?��*n���#qL�y�8l�T��P�4wd���$1'�=D�U�$�k1��T}K��D�Z|��@��ٶ��2�ͪ o=;�%��kօ��������&��ӆ�qe�F/��iO����`�XXy�r�����7��]��eC(t����.H?S�m��gD]+F���#�O���B i���
�i�T���v#�ؗ�Be:�����6����Wy�h�V��n����5���F�MΚ���$=T8�E(Y9���SS<�%D2d�����`�p��y����^fY�C�k�a�l�&t6��h�J���)�	�+�k����o`�Ğ[DY�->x�q�e�K`�i�i�C��G�J�,�ZfX��!�,�Z�8ݖ(<�;�xr�	��	�^�)_������A��L>��Ռ<���|�l��ըҎ�Hc����	)���+��q�g�N'�r�
W��Fd��Y^ER�]4YP�"�+��7����������6m �)���ٙ3�.����h���r@v\."	��Ym���5��Z�h� ��E���-���(פ3����ʨ�>� K�9$�afd��e�kA�����F���E�7�]t)�O����J2k��&П�Mk!��V�o��=7��x鬦������n8[f<�D;�hĜ��$���$����^�tl�W8�卛o.С�/�N� 0\g��t����h�k���4���K9�PCͳ�2!�ۧj3����D�Dr�3p~,|J�
��_J�?��P�3|��ˢ\��;CB�	��g�i���u�{"b%��5��#Z!#�u�:�iY��_(���;n����3�������es�[����X*��Lإ�L�s���㴋ጐ�	�֑K���k���@�(���V�W���s+��F�BkS( 	^���5�{��z���7�!��{�\�������)�,;����u�b��.P8L!}l�j�C��(��� ����#5%�-�}eA�x$kD�;���x�e���)�OC���Yp��GI�$J�~�R�P.�lV��%�,�\gIk��3��GM!|jc[�ۄd*D�Z*×�Q}3����FS�h��>�B)��+�^� 6�-O���.�������ԄTm�`2g]w4�� Pd(��h��j���s��.qK���xKk���dT����[+Lt�d�	ũܥ��q�,�g������0V�
a���p4�I֑X6�0ƪ�t$�wp�t��.�n�����ӌp�ک�o�g��z�C����$"�-��%�r�z?�k����jx��+L�������m&��8�18 1g��!}maE����{�>��.���ASDq�d�����%�Ժ�C�����k�y���H��Q�F-���c��=�A7��*`���K�H됮�hD�U��,r�>��&��sn��y��$6�� }l=F�IC�8o��Z���¾@���}�S�]����8�9Z��W��4���~ХP�ғ��ڎB�K3���e�i��'J٭�ܝk3�ud��s[�$�`#��o����b4�R���A=���q���9�[/�k�J��8R����:��I<H�3�TD�q|��/S��~j8Y���U�\�|$Zɣ��
]�IM7<\�܉����7�(|�l�{���JE]�\�Q&h#[+�Vn��ݥ3��`"��_W_
�Zŕ����] H��s���O\q� �}��}eU3|�<��*��|�q2	h.QQ��P���X��b����=�y�`���i�_\=-�Un��J��s�RM����bC9�d�m�S�o���;�����M�o论2Ae(A�������.T��X.�lȇG�uU�e�V:~mO��^Z�~4�Sʊg���G�����r���x}&�N��-rk�[��!�Z��̂]蛢S!��t	{ks��{d�4&����M�z���&jX��Cj�O�8oy@��p��8a4Hh"�-�Q�$^욮��&y��6��MD+��J��]���k�+�����(W@������V�+v$-O��f�Nf�@�&�(O���%D��
�7����1l�N��=��(b����0<.�_��*�G媵v��rZ��4�I�~u����"�~à՟��s�K�8!�LI��b������`��nl��S�擽`������K�Sub�N�zgu�t���a�dIM�k�t�*��4��#�)箞B�ukE�bAU���a�Me��|�$<9|�h���g�� 
D�IVY�w��Tݨ��LW�#�^(j�-�_��.e{P�k�F��4/s�'����l�_��)[)�H��,�\�G��X6�r��V7����;�P��^b<]���j,B��pdc{�v&j������Q��5��� �\O@�@��1eOr�r�Ej��b�}s����K�K��76�|C��Z��<L�~��G��'��âaXx�<�|�z��g�����CN�6�� *�S��ܭ��r�S���/���W�̉;J6��]Z`�="nqN��ޑ���c�k!��}\��L�D����p���h�˅ћءޚ����?�W�l�Gcu��Y����YWTw�"�.��M}�2:Er������D��n!#jk���X�c �N>�LX�OgvbK%��������;v?�=iC#/i���Ufå���Q|�,j����вJ8�YUvfӡ�����^۽%]I�,n��i�(ӦhN�D�\�h���P��9��m��Dn�]���� hjٍ��f^ˏ�#g�:P��B��|��va��?�3���I���oG�nD{�rVsa����8����H���{�=9�d϶���&�]L��y���GV-��J���z�<�'7/�*7%p�;�M��L��)�%���bk~� RT�K�-u5F˳��%��/���Gy��/'E#Y����?]Kd��U�zz�ǷO1ި�s@ѾP��1��϶�W4^i�mm������M	���s��a�	�QI�a�� _�`�fc��bA��B���_
`D���0���o�3}��cxfL������l1�X8ZH@�$չ{��H������+�Λ�iݜݩ�v���QPF}�.<6���Z�3��Nl�EFķ 2�6��zT9�[ 8�D��*닦�-9U0AQ��P��D������$�Æ�V�2��O(���� �|�ح3>i؇�*������d�yQ~h)֎�#��
n��Eqk<�a�o��K�q����c�i��L��r'@pǺ�����4$9+��,x��qz�����}�.z�z�Uw���;�?<�>�(�^�L�#?�{h�����g��$�+N
x�<�M��*��`T֟&v~�t������<.����gd�p\��w
*OLtt)P��jL�䳀�>��ء�{���B@�n��pmu�"�_�+�6ɑ�S�4��{˩sғ 1PL�� X�X��i���i0�P%d5]��� 'b#�́?׊��?�hVC�Ť�;6����������8��5��h/+�7�t_߻h��=�����+�ڗG8��=
F<`C�8�YT��"]���H#�)%jJn>���E�	fYy����O5Ѝn��q�Q��E�[�#9N��T[F9ާ�]��Y�]\��]֙נ�Lu���ܔ���{�L�$��ު���-�1-�T���4J��Ӟ|N�W|�h��R�7�j��E�Q^�L�[��JM��I:�	#�VU�7b��<�%ס�_����gQ��
����TڗT�v{�H�8���9>��*�Ҭ�xyU!4�[b�/dT ���;�wߍ:�%���~_�j09q��|��]��
��nt�`H��K��d��u]4\Dv��N�7�-�W�%+G|V��Ϟ?�(�Ys<8�֌s�L���GE���d5�]�6lMp}����4����;\h������w�<~In"�&���T�e<�v_��j����r���8�{��I:XI��S�DA@Wjs���o3^ӸM_Q��X�.��G��nz^��K� �kX}y�-����r���r�4m*ׁc���<�c�ȍMό������+b�N6!�
l)t�9�"ga��L�6SQ�.ދ�q<����='֗���Z�^�ߖA�P,��kx,-%.\��$w*�.f�T�)hwgR9B�h���W�{��D�bb�քDL+���p����vs��nښ4������ԏH��!V>��[Sɶʳ_�#7Do~�Yja���L{Ԟ�RqvG���Ǘ;�o�u���|ꭠb\�܌��j�����Q ���,-N���(���a������=���`A�e���Z��Z+��I8gvR�8��ĭc��d�_s5j����WGoҵik�b񇆃~
�y���̖u�Ò�G�-��m�'������̤Q-��_w�Ѕ�Cj���Ict8�r�W�'1F�%WY�i%緣��!���OPf�wԑS?�M(R�
Z=�]kAS~{ٓ�wN���U�lS��k�� ��2�3{v�^&'pŋC�iPHre� f�������;=<4��
'���]�-����w-VJ�������~��q�B���u�������_k$^!	ɀd:=+��+�r�h��(��E��EbW��Ư������~���cϓz�q�*X*�솠z���V�7��3J@3�h1h�����(o�#�y4sü�	1a!���l{�H����h����eO,H�m�3_���'�u]�ϽKŏ�%�	�q�v�&20A5J©#�����pB�@�ϩ�JX���2��������J�dv��{��� ��Cm`X�Xr��Z��S�g�lj�_��֖�2��=��q*��H�_̢$�9��t���.�5p���"�}�P�,����{�EW�#,m��U�Z���[)�зP�j���;����� ��uW�������M�F��9=gT�v�H	永 �����=I�����aظ|�4[8��O�1��.rޒ�40���0X�M�1[j���;��4=5~�a�CMu��(��L5���C���
E͝~�g/�%�ȁ�pS&{֋�;�M�8?���t�W�M���ym�:�\��DO�i#��#)j��r�Ч7�K����z��|k�4����#��6/��2A���j��/J}	m@���^�aGk�����j��~f�A���-�'(�G!iic����"�
r�2ߝ��np�hg��4t�-�T�&f�sܞ�?��3������0ڎ�5���� #�/`R��V*�m�f�HF��i���V��M�ͅ��W�:����0�;��ƻ)��T����5��
��H92�9���r{���z�ԋ��&���K�Է9��v�?c`�J�_�[<�]�g�)u/�����kb��r��T`�vd D-~*/ S|��(�(M��3[����T����{J��(0R�6�����9����'v�����u8��9}����P�x��f�Rq$�-�����#�Z�c��\o�����/��&���[3ޖ�At�HE{�G2N�)��\��	�=�4(���Y��Fv�~�SU�t�-Pr�t�f����,�wl�+@�G�{�{T������A�]�@��w���u������s��tz����.���ē�C-�s2�,�U��(_[Že�霟[�D��WYNS�i�Y�g�(]]�bj8	�������[��Ԝ ����lmB%j��L��3E�@��[���9����qԋ��x�� �;^�|�k�O���,�O�4 �r�ϩ�g٩�����D�l&o�-,���;�p��̂����1�����4�-v
+V5`M���b��l�2pF[q(�z�28_��>�>�6+f���]�U,�f �&�΃*�bx}1ޞr��dZwi���g4X��\M�h<�o�%�p�.�|�g3�I)]c;{7������M6��ije�����H�bǼjT��e�����ã:�nT�.u�����<�v��cфV����km�c�˶�k���_ڼ�kc���z8⿯��Ȓ5?�nRg����ȵ��vLsx�G���R2f������l#��,�f�����M#������#����>U��6�w6:އss�o���>��`kJ�y���'I�=%��Ee��w�����]˶Jt�@W�;hq��8j�
����j ��0���+�@��>bt3 s�˿��p�ݪ�@rbݗ3�Ʒ�b;���JjB�������
.�De��9S=�F5^R�#�1�Z3��J�z�b��� /�Lt^�N |_8�'W���`�r$^��x(�Dm�>��4�X��yi��&pPI��fB��T�~����8�������<��Ⱥ�z���E�ȶ����r��ӟ�t��31^��u�Af<l֜OJ�g_���(`��N�Ԃ� ��`,��#Aޟ���E�Zae���C��;~ݡ�ڱ?ʴ����>��kZ��M�J/% �W�ŀ��+Z��V�j��q��ig�T�w-��B�Q��>D|���4?=/D	���^�	�����B�Y%{~-6£O��`�˱1�h-7-�y���T�;д�ޛ��7�쨎�����b��k@�*֍�]�nB�T��d�kʮ}��W0�޹�H<�`+�d����@��c��
z�?��X.��w4�`,��*��V&N�m�c�*g��
���u���֋�ہU�P�[��$��H��vN�i��SsJ;���~�ӌ�_z��+�l�(�y\42�&G=K�� l�����h4hU�^�֦Or�vxٍI��4�iApre,&� �&Ws����h,�>��QN��ܖ0:`>v�8�6}��������a9�Ф���_0������&���$ �	��0��o�����ɔPv�Η���J��a:� ����K�j�2FÌ
�|5��%�7�}����2�n��C�����C�l�G�fOӤ�tz�X�`��r���7]��v�6��z|wm ���E�*�Y���dNk��q�rI�x�z�{h���uV�ƶ�>�"���n�3"� ɤ� �$[(O�Ɋ��B1/q��Ij<!�`����e2h�V�g���b��#,�?���7�����nd�e��3�	%�3���k���3�Rй��cwС��D7���r��O��Qx9�d���(Z+�� U�S&E8Ml��D�n��v��q����jegT4���v f���[�|%,�G��ˤF���m���M�g=�䗷�6��5�C6UM�r�O�P�������˾Z�T"S����#�ڞ\X��[�U��Qnv��pk^�ND�i$�E��%�|������3�sH�]�S�C��FS�	q,7�ŅbV�MI(3��g����������������T��J!p3=�g�W?�G�꽱�lZ�PA����J�<fL�����J�O�����6�yBU��)k6�u|ʓ���{;�o�3���p�#U:�lk�ɩrz���b�h���
��"�ߣ�P�4��q����A��V1XT�F��U�\�Wĵ%j���+s�L�;=�B���^G�S�Y��I:X�=9e�F�"`Q�)b�"�&1?���~���2�@i�ǵ�����´� }\��닉�%w �S���Ev���Q��	�<�8�խ�f��fu���`�Z�l^��I��f>�ҕn}EB�T׹���7�J�o�7R�7�����h��*)-�.��pDdǰXY�zl���
�E���|OIωǞ��?F
I��sU�K�?0�ڸ�b:�o�r�i��^���w�]Sq8�o�1�%�%0���FJ)&�'�)���u�H������*)ߙ�7+�.�y�LV�t]�wؕ�v�wp�">Y_wKŝu:{ÐI�X-i�
�΃�?<?�;3V]�h���,~H�>�+�'b|�Yg7�؍jt^�>B�Eā�r�_��l����U�8�h�<��]�3UtZ5IOڞ�oH��f�p��d�[�H�N�)�[D�o�����b�{�6����2/��;>5��Su��a5]�ۀ��%�񂚣'�����:��� ���d�>��v5?�y\r��6���e>&.˔4�j�žw�i	����?D������� hY�Z����BtXl@՛�M��8/����H���h���[6�~���u���kL��8^����݈�FG�$.�䜄���4�[��?Rܭ�]�6+?����S�$#,�1���j C�c7὎i��ƚ���Cl��M��.��L�I�R�����d��������N���	,zN���+�Q��Դw���O��g�t\ �0�l=�C܊�?ao�<�!/�O�������M�LW��<��>p0!�dS)&�������BJ��=�s�_�����$�I�Ê���q�;,��W�!Q��Z��~=�=��ټ��ϋ�nyF��R�<�߂��޺�]�y�r����^�.8�	ZT���MdJ-�m�6�b��0�����������8d�+�Q�d�":��]���I���(�:���x��_������r�[�	��*����Uz������� �L}�\�!�phTzdja��gWWZ�����L�Q�?�o�C�Zwo-�'U�Gh�P�����돼�p�Iٷ�Nw�Ct�<ؒ`8�Aht� �����h�R?\;�'����_����]A�4O�&���\b`e"IL�a"����� T�)��C.�cPmt��[��\�zr�Pc�F����!�e�՚^!���@,W��7����,�l��{�3vY�P	b�ce�5�A�I���pv���8��}�t����b:���U*6�.?՚-I�4Ƙ���J'??�6d�OX|-:�-V��=��3��z��:�)ap��|�9|�t�ɩmV��s�q�]#�qW����#*Hך����eb�i%��9t��#��?�)^Xx�Nl�юQn���-!|S:xr,%�kI�v�)�t<��U�����u�)7Q�Ȭ��s�9;�.�������-�{g��_~B�ve�ƽ�Yc��4=5�P�$Q��[9�j}���E��Z��;˲TO�mk�Gr�Bٌ��$��*�+-����wOs��f��2w�{����3h�azG���FJ��K���ư��WaKH�W�f!v��+W�����x8���Yi����@Q��K�J0i��_u'��t&яԄ2�����L��T}��/�\�Y1�7�(0�6\��O6�o5o�����5�A�K�jAg�éT�S
��X���%2s�賗�ح&त¤�yT;��R,;�Œ�).���]�l�
\�XA&�T�hX|�:��,�8!�D����)�1�����5Ʈ}��*&�oUK������k�}6�s`�G�F�kF٘�e�K�pv@�a`��z��c�L�1����u�e�]6���A�o8=�ܹy���JB2^[C�D�%��+�8�Ob�;Elǭc�3!aõP�yZZ�2j�+a3Ga>-�b�Ͷ���G��;����R����ɪ-�F���_r��,�ds��{leXI?B��y��ɬ�5��u���$��α6T�sӨ���D��t�|%�����u�ca�cYZ��#�E9�ٱho�W<�����PZ��'�]؝�N�j�1��t�*�bU���=Ε�,Р��S�2�
5j5�e�:���{5����l��[�=�?
._29 ����g��'�(q���a-�x�M���8�U9Ӈw	� �e�����;�a�~TU�.��8V1�	ͼ�d�%��z_|2�C���D�"	hj�(?,�b�B�+C{P�h�((������<�*u�CP��Oq�ʥo�GF�~�fl-e>q^��(���8��4��2A��P�����Ƥ��?Z��g�O��dW "�L�aIE����bM=�Y#Nj`�E���,��A���CPG��I�f�O�7�׍ŏ�%A�=����W!�q*ğ0���5%5%��P��w�����A�z�hlZ�mk��RK��, ����<��q�cQM�)�m�aH8|ٚ�v^AÃA������;!-CD]qe��z8W��>U�-�
[�٧S�ƕG'Ӽ����|[#ð�YTg��X\*�o�Fvʄ�1�NO�9*�\qrZW[�c����8ӫ.��zp�8
�Bkߨr�#Oe�~L�A����Tb4򇽫��t�A�d/w�(����S�B��o5��+���=���0�Ҕ������5���������ʝ`m���y��O�'&k9�ފ�I��>�{�O�m>FB����u9'!��?��7�+�"L�F��"6G�>W"����q7!F�l�U������X�P��_FS�#���� �>E������Du�]�K3=E�}+�.�;��LI��n�p�>�u0�ۥ�/�]f=�޿�W�?�iv-O����*��5�mϘ��)���d���8�WKdp,f/�˨��~
$����[+�C|{��_?��6O��Q��7
�XB���'ܛ�n�+��UI��"&���"fv.	��f�?���&��D	�yzr���0&{G�[G��2��G ea}k�}&Pj\��k��oWI��}r�u����[¨f�e1A�嫨���Αja�F��E�a�G�����]�l�����w��-ů�j��6p�����n,�n����{�2�ܫF�P�4�֊�>o�{�cG�h|�I��*������(7�78C=�Ma<7��
1��9�o��P�.���d���hw󕪃E�)�P����T�ϴ߂�︔(����eBN��0�ET�ԉ�ȥ3�� ���fx��ë�2!/���F�F��mP�%�nL�s�|,�P	P ^��s����=���q| vؗ_�f7�|}DI���XVL��b��\PЮ�ꭿ\ed�T�=���-*����N:���z*�N�2�ޞ��1G�0��˫_��WZ�͜S�^�	H��KN/ieE�"ƽzg�k�?�����S t�@�HL��n��I�kD�mM��9r:���a�Ip!1���*^�}d�PW���<�G�+�Y��r>�Q�ⱚm��PD�;�Tf��-��-��U{���j���?ֲw���$C4�]�g�4_�p4�v��d��H�ڣ�����g��>&�4Ԭ�E7�X|A�8�0���+)�ܻ^�0MG2���[��/�$�ke\ZN��5��?�`�D*,�|�	�'�=7�'��������X;F�w���p���_}�y�}rO�jE:/�7�t9�h0�:?���9^�8�?r<W������Y�
�|�����][��B\KTY�/|�e^s?>�{������K<!�͛"o8��Y��I�I^P+�4m�vqFM㏈
/�SoL;>���:$����v���S�����}��V9d�O�Ѥ�_Rl��� �z�\�Q�=��z#p��ï�O$��j<i��b(���sz༴��d�V�f�V�rvu��׎���R˃�ӱ��n;�e/MZ��
�� ��U�~�a��Vd��Y��xy;-�j�Q"�ږ�8?�gkr�[!%W�����,�E�h�����;��"c �y�x�X0"�?�Al��#����5f�6��2�H!���Ҙo9>�}��Q�d����\-Q�9R��jE�X��XT����u�/s�X�����JXX�0?���14��],`Elh��{:B�|�V4]�;ߞ$�A��VWz7Lp�㪆�Q�|������h��Al��J91�I;�Ĕ��6Lbu���e���'̢�+%��E�ō^Mt؇&�H�,pj;��v(}Wj.䔪����H>���cG�i��'�y���r�1�4���n�����l9��6�Iy��ߑ��/���痔T>���v�	�����P������(���e��@2�-9�#oT�z`��y]R͋#]��_@�Pí��[D��� �f��F ���T��ghO�M^$ӷ
���L��i���	ž�����������z%'�����C� ?�Q*�����8��*��۳bK�=���⥰�+)�7�ǳx��4����M���j�0��j��g�b�Q3���o]�Z-".�:c~lx�U�G��b�	A�zb��E
8�cn��_�%�2���d:`��=i(���w��ۨ��za�ߑzZ��� �@���L�䷫,z�� �%�ʥ5��J�IN&�8��O�:D��./I��6!q?,�GZ_3[�4Ej���p�ī�רf���_=�J�P;��󁸙=P+��kS\0k;1�g߿}�����I!L��횚c9���},Qr?6[���E�՛x � a��x�"�o|��k��Б�y�Rn�C��*�V_ ���H.�=�G`%nJ�D�mG�2�d%PGJ��&"�_�~�f��&)���3��"Ϋ�"ё�$Amg?�����&����VxL�Hʖ	@���`�l����2,���+r����J�e��:���=��z!��O'ȧ'ToM�!l����y>#���@'֘7�:���1�͈qaX!E���#SO��A����s�ضtX3��gh����yЏ;Gi^:���>��s�h��\�Sr�bUF� ��	m}�mD�h�G��T��\��|ݥ=�Q���o�������M_wl���e-��U,P�M��1+vQ�c��ᤛ��]�c$�J�#�{E^s~Iϔ���������2�6�A��^k\����LBq�cg��\��s���S��{�
�{�+�/�Z[�E/�#��D:s韛�h�l	6�i�,Zl�n.+H��w)��q;h ��~VLA��tZ�囏z�;K2������
Z��M$%7�s��aiL��~E�/�������NÎχ'�Qʨ��e�x���j���C��ؐ�0��I��]�*پRa��q���R^0����f�V�,4\���y� I`�U٠�D0��*��$��Wq��� �:�rV>�f�~����,8���x����Ng�B�zwN�5N���#J������y�����;�������;~B¥�˚~lɸ�̬�EH>����L�|z�#��
���	5��e�Qi?7I�;$�?	�_���}��nO
"���7�^�$W�V��Qu��r����c	ε�o��a�{"b�:Ӕ�:����K\eȒ�5�%�#�Vc��5K�B�8(���y����>��J����9�ځY�Ј\�s���Vo>-:��� �pmq��ta�c�BVu7x�Y�Vu��i�kb��w�y^*8�_�6�P+��
x 5���8����H��s�����'GR/;��&��W�r�W8ײ$5�B��s#G$�2���oz�i����v��Q�0���32��%��M���NX1�f��.�����cc�����PwBrv:�-K^"�sQ37\�W^�9-u
=z�ȸ�7r���/�9��'o⃘)K_���w���S�Qˇ3�ֺ�t:�$���1'����Kv�B����G<BEKN�4p���PlI���!�H�y��W�3I��0���4x��Z��1��r�풧@j1�X�4��
�2�mG��)�f��d]`�K��R�fL�U�Y�)��@��c� M���׬�t`Rth졈�1�L	�wh�^/y�;T��N1��_~�)�ǋI�O>�����Ugߒ����C���ݔȓFة��r�ѐf�pԦ2�P�3��*����<
	]�(ۍuzf�@I�<�j�~ܙiL�^��qIY�\ [�ё�9�	agr�j�铲��,���Ȣ��� ��6��dz=�'�p�q8�C?}�s��q*���-�Ey�(vI��i�G��Z$N�$X˝��w�=��g��ܲ�݋�R�����єe7�á�J�����{rBJ�&ZpAzb�F�UUqQ�q���Q��(W��*Mt�ݾ� ��>PؚP]����[�}@�sw8��jiq=щ���_6-c�g�U�Lv���A�=Y��Ԗk�w�����^���'��5Y�!��O��Z�x̃-�Ѷ��{r�y"�-�2�Z����u�¤��@&�n�5��G�4pE��ع	4�$�#>�I� �ņ�����+"'�1L<X3�͡��������E"�!n�3�vyq���g�ћ�v��6��$y��:h�JSsP��R�}��{�X����l�����!�`ZRAW���
k�$�|�8���/���ڄ��lAL�� ���%�<���������qӌ�O�0ܙ�m7O�W�g}`��Nq������2�&�;" ְSdLK���k�nj��'l!\�d�8G��HL*�21NN�gm���oln� ��*.�'t��9	��|��$�E��1�^��[��(�I~Y|!d����k�5"k�f�0޼�a�O^TX���x���L��^�����n�p�@�6�PJx��@�ա��Ϝ/o ����v�Z@Z����I�x�,A�!���W�A��*�ۘ�GS6��:�/��B=N��
eR�ߌϪ�r\q\RM\8<�.�X�^�E:�e��j��#��t=�D�|ɖ�&��{��eM��l�S��p�Oi��J_G���Lf����u
]��v�*���юU>���ߓ�����o��?ƘAPQ��0�#2���e�bD0�)Fl���E�-2f-�#ve/a������!�����k�<yZ[^m���_��g�:�6x/��;>B��Us��w�3�	rQQs��)�|�s���	��f��)�p�a^�8M�b���=Ɍ�P?;a2�[X�q�7kd��+R�Ԝ,�U��C-Ւ�T�a�7xƮ-�B��7k����[#2���$wG'�7'�-S�|��g�(L��O�|��W�M��̻��CW/y��Hgl��n�F]d�X0CH�o�;~�;*�h�C�I�~=�=4;�}qHu��@(X��^��)"�T�I��.��HG�nT�>�~�U �a��9؅R�J��:��Q�[ب�?Z:fR��
�b�5/��x]�)��3[<�vl�� �"�	�A�П�A���Vz��cR��c���H���B7�ck�w����F��Y�m/�=�茏^��V������cB<���3��P�ٷ�UPY0�o�i�װ%=���!Y�U�%Wp
�C#
bwn�j;a-8IZ�Q��R��{=��=�)�g�y�6�a��u�M�#D�{�m5���O�����jI�Z���Q|L(�`�ʝ�U�jS'}�F��$A��H1eT��k#0pl�%M�w�3s���x8�OrD|�xV�^<<�ϻ��Lچ�u4�������:B�e� Τ�l�����p����/�$����R�C�
�b!�t���ph���3kΤC�O��f!�O���c���,��P ����Z���a���4��W���(����'��5���ym�1��4!��N��Nj�n��;�����.,/ x4g��=�-�9�x揩.��J�ܢ�~���$	C䫘v�չG��!�%�9(Q�_��?v~|J�ص's撥He\H��#
����8W�0�!��
߄�Z[���q�^��h!�%i"�B����e�"d��UF�I02�	���;~lK!��Y���H_k�e����Q��N�	���1�Tn"��nEgl
�PM��,��A'�잒�K`Pc����d�U3�_���nHwV���e�J�.{�<v��|���{�,��% �[0�'� ��a¥:
4��L����V[z��ڮ�4���V�q��!���u65�w~G%����!�Ku�����ȫg?���7_ `����U6���̭=�d�z��a��D�O)wt�jH'��b��wK�� A�E��<1�7&�D%]�ݢ�� ?m���8[��pS�4��f����Elİ�;]�60Ǿ!�ʧ���}_��6�� Z�r���������b����q��(ʈR2xA:��.�^l徳0
�Q��˞U�-��+�6tû������r=i��F�/3�F���?~��ӏ�sX���f��SAЯ[�"�(3$?�+�aC�)♕W��Q���l[hVK*�4��N�z	�l�ܠ�iD��@�Y-����	�i��m���,u>q����D��~���u�����M�q��<�L@�7�^�K{��+� .�w� �F��0-#ٚU��ʛ���2���
1&`�1*B���߿4�Xj�_;�
L>���]�x�S���!p_�Y�۰�?HuF󠿌�:��3�}tpH�\t��,�� kG77E��S|z�k-$8��p� q�E���ϟP�v� C�8�Į����S��qj �t:%�hwEfFc�&���8E�����u�D���&�\f���f:�3��֎��j���<U2�3�;;ƦG��sw�K�I=�(
F� �%�5z����3�}��I���y:��	T��1�#��l[}Gb/o��Ԩ}��2?g&��Ke�L���U�輦T�t4��B�0% ��g:L��[$!Kv����Bd�,#��
�}Ȣ#����-�b�cDS4#���/���~)���p�~�J̛�#;�į�ݙ�T%b��D��y��y�5�֐6����K\��aa�N�כ0q0���*W��8���2�[j���ēS��F6sN�|}vr���#K�MM⣼�2�V�*ɰ�٫��?�$����:TP�a�*�k���2[�����q�mŁ��e����w�`dI��w� �2sq��Ʒ�}v3�b�'i�F�!!�}#�7N<tjq����=�w�{)�=(��������b�f���Y��r�8�G��:���[h��#@�òq��Ŕ4�ڼ�E�t��U,!W���o��w("��ނoB]�\v�!���� �CR<@$����|��R%�u��K~B힌��ܓ��!��ߪ��wj�`�G��c>�2 �����Ũ`�H� ?w: ��0'�BL�R*�~yJV���O�1I��SD4�(�z�Ӑu�J#����t)Ɏ�;���c�O��HsF{�(��RqR�"�Wvo�<���L6�sj�T��0��.)����)�J�Mr�m=�2YJ�
�jK�Z��A��R�N+���f�TϬf��{Vġ9�3�͠b�0��_o�f���u�{����`���2F,�9���V2)aOq��e�T��M_�.I����i�Jzqӏ�5SR^��g�<�r�!	��ʤ0�J�u�,������1֫���{�i�U����S�PǴ�x7g�0�+H��+��o��h�Z^ġN������l�h$Mq�a����T��۬�*W��=���4�]�&�=�V:%Lu#�ך�H ZɲWPuM"��?WqBC����w�|p֠1�؃l>簕�}sC�K�~	!�*��`E�K�h~���Lw�����JT��_/Z�v��6�_Y<�2_�ӿaHy�V�����Q����h�/Y�
��웧/��`.�L�!�~��*,�;F�	an!1�mҰ�i���jݓ5��;h��{�v&��B������Ah�qp��ߝ"q��Sw�6i�Tr��Y���F�8��7�Gf�/{8��b������FҮ��x3��`;i-�Ӡ`�C�(p��� ?�|	CLv���ז��kk���c�%� �Us@�X9ȕ{h����72��9ѱ5�M)��^��f;���·���*����&�О�����C�v�ad��_�����A�=�4,*���2d��m��.oN�R#ޖ�8Zz�wz�[6���ɇ{E�� �v���#t��:u)nP��d��3]V+U��!�Ն�{�K?NrE��l�����[P��-V�+�Z�Đ"-����D�Lw���C�S>�e��,
l��$n�q�|�iIi~�'z����m�hz���i5��YA���T����i)�5R!����(��$��[�D�esT��%��B%P�?ɤ��E�A��7^�S>�d]�Ȇ��i�}׮eF�ͦh���wC""tK\k�u�5}�s�>4L�W稤0JZ�@P���������>��D�����Q���:f�X �`�$,���WH�17�e�#��R�5
���6�:�V�[,���Odڦe<<����Қ��5��Q���E���}S���<�j�,攟�? xϯm-a�ΣjE��1ˬ8ő�z��~0P�k���4i<��,�Y'-x#|c�(?����F� ��/���^.�-�U�͐�ۀ��G����yo������������ʍ����d̼����\P�AH�@�� ��$!�Ұ �|�(���H��_�Ȯ�ĳ��C�9M�9��,�F���"S'�貏����	�� �+cޛ��P��$���UAR��ӤW� M�˒�� �x�E�@��Ή+�
*��ޕ��m����Om�a�5���W�wרD`M�*�K��R�ȎL���EgW��W��r^/j۩��r��� `�����u����j���F��ŵ�*�Xvq3����#�M�\sQ�m�X�W��k;�R�	[��'�����*�X��b�b�z�"�m�k��{��q��6��H�6~}�GHSa�b[���L��W[�a�!�M��)�X�ê������j2��jm,TN&Zԭ���;6GM�53+��t�VǹN��&��#��[s'���Ks55��m�8��Y�������(�B��$n�Q� ��e<��iݼ�p[aϊ���f�]�H�]�`54�"�vI�����?��q!�Ѥ��T�V��]�!م*�r���\��#D�Fa��T�bK��f}Pg����"M�:q���yjw�V)����mY79sO��2�hn��0��ꋕ��
�(�L _��C������Mjh1ѕ5PPn*X���G�T\S��z�Տ{S4о�L����~6��%?0v\��j���}���Uf]�5�����dw���4(�E/��A�6k7@Hƈ-(?����3�O��\��)��Ik���I`ͯ�aϽՏ�.te�*�����F���1::7�(0UCì�tc��	�p����.��N�0���˟^.�l�mH���U&��,�����8��欜�S����GC[w��um��C��4h�ߜ>�Fx4q�X��V�Q�)����Qty�o� ��O��s�0�˻�~=~�;M'1���s�귓T�Vg!L����r�Wg��h�(���6�%�ӈ��aȭ��ɬNF^�mA�W]o��t��
��;1B�"�����ŚM{tG�OMm�$�0�������Lq4�s:�v���Z� Mr�HX����1����,��c�**hC�Nlҷ5����6T�Ը�[��������$�
28��_��RJ��k`)�m���IxcAi�9�l����or�����N��VWFL8˓�}�{����V�M�w��t�#jע2Dr��ky Gٔ�]
��E�h�p��<0���1#c,2A�{{���h���<�B�nDQ5nJ.I�|ttТ���M-��R�@�U���%]�	�������c|�?_�.���Q9�A�T�~p��ۄ�C2�BP��3lh�o�?K��`p9�B�l�6=�yht��E�-i�ߠ2>��>���I��z�mA*�h&~z6L�н�����{�1��B��m�X�
� ��G�`�.5]�^8�B��PI�]G��B��x��|�nI=P��W���l�Z�BN�j��[Q4aݪ����Ґ �n��������J��[����J\G��NZc$�(���c�F�u��{6<�,p
����$�Ad1����	���Q�r�6"�UM`UR�恺T���L�c��T����Zc,%��2'�<U�t��8��7�x�n�~Ī��_<� b�$��}������� ���Y~4�B-�,xSEz܄�܏��U�ݷ}�Em�4��4?	8�Y��B&��̇�-��/�>��[��A��(�NӁ,����Qt��.&��p���LI�V�����d�qf�Da{F�3��ҥ�q�n�gٰ�T�`	��Ȑ�{t�݆�m.ˠ;�F�!�薾}��G�`u����;����~��,�����(r�A��U����XE�E_��6m��*`M+�h)��7�SSY7�������dA<�U�wG��im�0�u%G݁��3�Z�v��m\���������s
޲�	�?�5F])
pE���""��h�/��|INϥ+m+Mp�Y��J��`�T����'��t�=�_�9m����˃'U|,= ={[��m �T�2p�9��ݸ�&?6tO,+����W���ےti_`8��R=�.���ڼ�gkP�"N�N ��>�1d���aĄ2@K�ͬgW鵆�[�z��hwK�r�~}������f[Z{����>�X����l�Y�	g�j�f�<�iTԞ+����/�a�`]�Z[oI�z���#����m�)N˨�����:`�o��+1+��_ʘ�ۆJ6� �,ơ-S�G{${xr�����/<��:���(��ۢ���7���ש���+��c�$�J+{̠������~6_w��%XT&�=h �c�~�.��ns�ɫ ��9�(�p�/4Z~�>Op�;88���Z���ia�ۙ��7a�m����Z��W��=�4A�X��������ϟϝ�3�W����VF?��P	GJ�,��l�oW2��Q���F�d�+p�In�.�È[)���Ԛ-��ܛg3�iHC�|�Xys���_��~�{��ߊjO��Մ1��.�g;�q���?f!�@;q���);h�����(ryRվ���;`͝q�f��*zl �kGe���v�܉Ky ���� �Dy�_���>�ۘ(\�X��~�'�����=o�e�����K1���\Ut��~�zv0��T�C�zO���\��f�Gw�����_B�����Z���J�V~O��|��聱-����H+t��$.dE��|SZ�"�1ϲL=�5��_�7N���_�8�S��q�A<�	Q!� �`3�P�[�Z��~5ۆ���ҏh��;�n��h*��ڻ�%���؟�!��%'B}�Ǔx�b��?JU��$6|�t�cڈF�a
��t��^4$h�'A9iư�r͞{�����<9.C�fUꀅ�)D��uK|��v��zܑ���q��ON�0����8��_X�bs��Z$�� �O����T�|_ʠ��&}�d�w�r�O����l_T[��|���<���>�#O7�?�+����1��p�j��-0�*�����{Cx�ܖP ��~^��l�ӛ�#V
ގ7h��ѐ��������(����E��Q�������[�����oDm�-���3b;0����L���mz�>V�
��Ж�}a	�z?�ru<�iY�4
�]�ւ�J k@c� � M�1�M˪'��o���)���v���Y���݁�E��R%)Eb��D]�����i1��w�s�/��L v>��@���<
b�Ϩ�l=2"`>)���I�������M~Ab�}2�o;5�Bt�#���h�R(�6�U�|�U^�\}nf�L��r��y�iI�2s����8�l�_0�a����*����'�u��k����7�=cǬ�#x���dx�]ǣӁ�6, �4n�
q����������*��i�:���U�]�����:)^W�	)S��_��'��C�R)��.?G�%���Ŕ�=8��Ͱ j'lu ˣk��\�m��'8$q���i��6;���F�'�
�'�3�:��8I��i�ϢI�}�eb��"u�E���D���M��^E�|�ѻ����;@Ee5;��a��W����'�������i����L���$g������cYf&~��,��3�s�=Ks�~3�酜�j\~������"��e�E^Ć��o,��)]+-��B�kSH^(�f��j�U��D�P���4���Ѻl�h��T���wc�_���/C�O.��eq���;�j���/ok����"� 
"O���t�F����g��k�"B�Ĕ�F�����$u[���1L�c���K6����`�y��_N��L�'՟ 9a�-���F/�r~�_Z�ZG�����{s�D��F�.�T2?���&�歩s�/>,"�����di�Cێ:�!f�nǍ��:>�j�M�ԗL�rR
X�����š�M��ʙۂ�-�Ţi��F,�m����;���r�M�t�ؿ}��?����-(2>K�@E�$Rrii�%1I��U"�Ğ�R|��;�?�:"Y@���}>���5>:6I�珒W��E����&Orv(����R�o�ߥ��Ⱥ�'u�����IՀ���MJ�w7~��|c�c���p���`�.����U��Q9R"zY��C4=��]�<k�|�h`�ډ���e�䁄p�g����)z{|��>u��X�i���Y�󱻑�I\�m��sx��٠�H`e�Qj>Ǆ\�4�i��8���:�v��1�=�y
��E�` n�^p�Sz�=�aJ�i��7�-���RI���
�ge��/k~6�U��eT^9?I�A������z��6�%+c���_l/7���?Ғ����+�s�O�R�{ݺ���3���J�hWH�����4�Q�wK�n�ObD	1'�s7�Xu|S��l?K�kWj�Gr��\I���n��e��Hg0B�<�*���fd.����r��s�,#}��>^^�;I�0�����a�����u��?[Q���F1Wg�������u�����ɓ���Ɲw��b���pi)�|-�`:�ǉ4�p���ekrU!�M=n���6!�S�z��X�	UyoLT�<�Y�����N���N�b2��[s�aGӰ���+W��z�4O�S0�M�Ƭ'�@�F�c�<�x�0��dɗ�܃��_�o���	��i��y>��H��})���u:�ͧ�%r�:�pg��w�g�{|�./��'Pƭvk���ИץU�Z�~�s-��\"�J_o(��zH�Q�ܔ��^{�԰?��<Q-r��4��J>0�_v�fQ+Q�v��+�-�b��IM�D�͋@ϱ��0��ɏ����h�6���:Aì[�]ʇ�+3a7�lѢXSk\|X?�o��)Ɓ ��%��=X��tF�4r���,��O��Ί��n4��A�͘b#�a;�~j"j%���x�D3��aҙm�G���u�ϓs�	��*P�Z�T2���R���@�D �x!?�;f�q�C��&��~�mT8���xY�}LIKȖ%Y���2��Fg҇��X���&���n�l0�z�D��xs����;m�h�ik���`	@%�ur��U����=$n+�}�4k{S�K�o����L��a���uA��<sE��{˵�����?U�1�3��5�էy��5�VѺ���︯�����}Zi��u��u${��3��عȼ�Yo��ӄ2@;�ʄ-�M��-�`��hǷ���ӷiJ�nc��+����*}���xEa�V5~y�٠�(���m�O�0gM�=2��z`1�vɇI���G�	�Jl/5�.���m��8�9ul?�����,�J!�#W�z_�vt���WQ��S���:��X�T�K�tVM?NO�K��,��򄎫��V�����B-L.�0Zp�h<�����*�`v��R$9)�}A�����:�lN����:J)�G�3iu0�d׬O�p�d�.z8@�
�yC6⑟|wvnޘ�t.4��`7}�rdwBzљ�'���ZU�\������挪�,�(緡a��t�R�|�¡'�*�)���q�T�:v�<Z���,���١P������`}�,��(��}��)���t�?Ji��1�č�#�FU,E�G��􉫝���h���MUؐ⑳L����d�b&Aޕ�x��ȵ;���s�ּ$�Σ�훅�υ�=����<E�]12���h�O*������j	�1��v��Or�A�BOW��7��B�}3>E�/:Cu�����l<�gfx�,�{I54$�©�F�����2��8)7��'�_/7|J>�'/���������J�6V�vh��Kj�c��/��ai�i�ġ7�v��8����n�0;�O?@m�6��?�3������|z��f}RDe|�M��J�t�����j�왩1!;%������8�"�'yZi��F�?Z�MQ]U�e|QB!��3=�l.IL\c��H�A�N����J���l2s<oս��ɽ�a����-R$�Eę@/h�~�i�ԃ�)��=�>���z���\��B��H�x�eL��?����{h�SW֜�������2�}mA�\;r�m��翲,Ԏ�Hp���+����ttJa�9H�m-xX���ٛ��)Sؔ �~D�(Sة��\O?[���[�.ߨ�=��ɠ�y��ڍQ�K� ���ܶ�v���ɰ<  ��!A��QB�#�%�K�S��޾ �(�m�H}9aڹ��k��"wqՖmL�	5��_#��Uu���z���I������0�d���l�+eI��� >�*{ƒz�3z��E�LҧGw���˗�}����!f;��;�W����|��'����ч�c�=A1�N*����ns�%�\���_��Fj���I����|@D7!ɶ�����<z���*� �����/b�i|���K����F������u�y�#j��\H��óp)x�6���.Ĉ��?Z�s9(�
�z��)���Q|̵����,$�������D=>\�9�é9ͩ4��N�)�^X�s�*G.Q�~�u:H���l5Mċp��,�F��ͥ���M1S�𩄯y�-E#o<�; �A��8=N�Q��bס�F��Q���X+���X7	ɡ̙���9U/��TYTS�U--c>5~���?�]��1�����M�]����KKԁ#߉*�>i�7A�p���1�c�z�Q�����6~��#g c�i�\��6�������If*A �Y��}�9P�HV�ʂuґW���
�n��ĳ��Y`z�E��cv�j�ܴ-Za��Ta�l֔��^�2e�/�,���GX��7b�:� �����lBz_d���&ž$&��V-�4����AB�dv�u&5��uv��}N5T4�an	B�*{(]n�;��4v��7�7�Z��}$A�O�8��=$.>Ӟ���qk�\xUJ�Y��bE���4�#6r��:Z�X�j�tF��$�3.C��@�À=�%#z��)R�VT�G>����w6�~�?h��A�Z�H�i��d�F��GSCJ��s�l����]1SuNQPN�C��' �5�O���_Њ`��Yjr���v�	�4�1Z/��a���ɐ57���F��_ �B��P��W i��g�7��/9���o=���.������̪�5�ܠ�)ᅧd��I���S߬?�l�A6q��}��T�<���4��&!f�쒱�2�W�I�k���)~B�7�˵ �o�}8�dt\��(�{��.��<|`�~1c�W��05�{��ݢ� y�J��=���1���rʋ��1�o/�뵻΋ Z*�wJK��K���c�*Tt�%�̬���M��1>��W�OO@� E"�럕� ��-���Qi���	�?�(h�V��7�OD��������*��uS�ۤ��a�r떴�\Jݒ�k��������eX�3�� �4T��d�7���t��J����`a����\����Ũ0P�A�8���+rς����|F��M�$���f���Nր/^	�f��i6.~&?!�
����5xxI��
<��'C��6�u%����d��"�t@ �E��y��Nn>�7���7/P$`z]!G�کN��a���w��ĺh�YCe���T�~o�C�{*�q'7	��K�cE�R��5�"p��j�f�P:==����Z���3J~Q����4�0�th�,GLY����ۼ:>|9p�S�Z�;���t�P��Iښ�HZ�46�=@���}��4���q�X)҂��$�FK�f�2���Ey	� U�8 �O֑�.���'�fͱm[~>ۜ+X�������GR����+֢���!	vÆEư������o<Z�e�4��|�|<gI�f�]�i;��|l�Y(:��w��'���,�}K�P�p��BuICe�и��'��H#	6�ճ�sc�<J�� �=��"G}�9MTZ�;<�D�ݦ��:��D�3u��ke��5f+x�fB�<V���e��}��&��枴(����&�h�Hˀ�0�Oo*(�+�A���x�VǑU�6o:v2�j�(|��kl�ʻ��܁Y�j��-+����}�U�_�F���i��L܎�Ӧ�u�gr��YW�qah�ׁ�V�9����7����U�]uy ���*9y� �;�o�!��)������SIگ�㮲o���CH�"!Uy�K^���MG��@���p�e 7�����3�m�����X��{�˙'HB��=O���ln�����=�Q�d���2��}Gvw�G��:.5�K@��м�7H��qZ�_ ���޴��KН?}p�p9�PT�PWA���斍���@8<���k��r^C�r�pK�	�Px���ߠHf�~� �:#��%%�JM=���W��5Zϵ�����_��<����w��f�����g�߅
ˋa��g�Wd��j2Ăs�;�7�6��t ��o:�y�E�a�M���:��ɘK��4�ŹrI&Z1r���,�M%J�eT��Pa�A���&��fk��=3�29���֛���/�Y#3��ݛ���6�h�:X!�_<���]e�z*���ھ�0�B|=�zw; �,ں`%���x`�4���M�jb��@���Y�T��?�Ԣ�)���.�zs�g��+��E�nB]��=���i��e�+̡�8�2����lUU�@��)�+��/c$�f�ltQ��^�����!�yK=D�="��?PX��*ͮ$1P���i��U�kG^�=8�qغ�����	��d�SS�-"��I^~�&0�~7���1
YBxj�V�<�0m����{�����Y���ڋ�RzAEUG��蛰����|t�N`B��j��T7���UG:��⇄_�M7��_��x��Sq��ٹ�>[�+',�I�w+q\ I��1�_�ƶ*���U�}:ڃd�<R%�`%'f���9��7��|���S��@��z?��Z�C�m���.�
��;�6(��p����,��n�!�� )M�yZ2��-�,w*)b$���[鱀���5��w�a��`!}ţHlm&�q�yR�%���F��t됧O������ɗ�*5�N�dds`uH�D���mg�j8�-��AB���z�'ib����b+2D��S�i�ڊ[ʸ��
�_�L��5y���NdQX�'T|r�P �T�|����_�$Z�VeǒtIٟ����na�����Ԡ.��Yk����5Yxw��^�zp��Z�`I�{�s���G����4i��`�}�$'�צCv��ve�qd�IOh���`y��J��9sk;�,9��c=���[�����ɘ��NeX;s��-c1��|��ڃ����.�]�Jb��&�kᶉ��,?q�pґ�E��U%���N�-T�JAI�`����$��WH�A�٢��Q
��g�RUI���+B��6$#�!3bsa��Ћp>E�!����#q/�_�Kqs��i�c^��pLy��;��ig���mz@���6Ǡ�~���4p�ߓ�Fb�9�	˂�%����̇�u�Y���_kȷ��,쎮:�*;+�O�Z��8!�r���zx|�ݏ^C�V���z-$���������V;�c?S�rW��*Ό�j�4K����F�%�}���:��4�ÌdK����y?��c7���̻^�Y�y��^��*�\�NAe0�.��(BE:B!3����v�E�]z��M�d�@TFP��%�ˇ�"��I]����=��>��z*��BC)D�"-t�3!:O'���6!���~&	'�az��P�O�%�L��d�i`�����m�܆�)w�R�Y$aW�y�+��#�(oh�ԛ4�e
���y�S���>s`i,�o��g~��ʡm�q2�z=�������ɋ�MZ@)��6&�6����2��6��qZ����U詗�AW��!�׋s�Ây������z�2�s�� qjudz������i5�P�*x.�w�%�����U�+r������q>�ъj�a��*��rĄ��qg@;��x�6Y�~��]�]���υܚvi�{4���!{�0��+�Ǿ�?^�6�{�U���p���$�5y+��c�Ҹ�7���Ɓ�_Y�y0ϳA�\`�:��qtP�膝\��2(B3�z������Y�@���&��֜;��FZ�[�Y��ֿN��q�f��ZA�NzU�D�Z��̲Ώ�p�����+<>;��m`e7G8:K�������(m�q��S��Fz��E�W]z���T��6e�S;+
V��I	fJ`����0n��D/��V^��TgU��	����5C�l&�uS�.m�,e�kh5�Xx$nS�b-�M�"Z�Kп0<����í`6��OJ�3��h��u�$��Ö����E>K��k3�"�
�w�Kf0��-�l��^�͏�����L_~�5�����f�@�{B�cm�x@UK�T�����Gx��_���SL��Z�L�Z}�6�q�PO~�t��&x��4��=KH�k=u 72�1��w@��nR�P�����B?�W�no[]<�H�ܛ�q����<r�l��uU��m�N�<����D,����d��s�}�q��%_�)��Z�n��̌N]]���G��F�r_=5ܪxzώzVG��c*���)�`��>D����'QX"t��Ű��m��`�[�1��d�����n����_�tO>���a~�w����
>{5伥�!�8Ń�_L}�X���t`�ߋk^Ĥ&����U˅���4�vWuz|W��-F�u�!��C{Y��7io���0�l�B�H
!,��� �N���[p%@Ij�F��n�H��)Ui�u�C-sZ����.+k�`f�S�s�s;���M���yH�IAh�\2�d\��������� ��i/�ȩEg�ME���6��k�U�u�2�]��'�h�v� M0��"�����Ƨj��h;��9���To6�3�ƕ݅��%�ym� WY&��Iމ�����#�##c�j��(��l1�Đ�����G?�����:mbL��\���2$s�Z�ţ��+Y1Rw���[�XH��E�Φf��+%���͖�i<��Y"�L��8���N�&�
�5p+���Xt�S��=:UE%���Uy��oP����//Q�q�O�вo��KGЃ���n6�.��S�Zǜ�y N�������-W7���ߏ�i�8j�o�����'��C�T�"h�k��Q���\�� �yhB��b��|tG&5�  �#%�H�ӏ���Q?�e�ӊL��h�ʌ��T����v������/d�Gk}��e}6c7�́��Ȥ������ϱ�T^n}UEez=<3[���)CN�1��u�.�D�YÈ��8���l�e
6����e�W�'�iV"z8C��m������k*�f ~4�������ˈn>p�vƬܵ�A�9��I��ُl>Ro�.���XG��~z�F��7�5~���	��z#t�XL	DF�_xڪR����lc�l3lv�xo^;E
說.�y���MB���:=�����_äF��#&�Uŵ�P�,J�]��;�*%��6KM�Z���E�5���
"�K�m]���P1p�bxY�o������{���w�f�s<��YY��i��k���M�ǧ+T��ez�73��r̞��z�17�����7&$U~�4_M����M!Z�ZB�/#���	�0W�x6�)�3_�������b�
�[f|lGa��>�iK�Q~��T5��آ�* y)bw�#�Q���f��E�����%i���h)���HH�&�A���Ј�'Ç�l���x�FTԀ�>»M4��y�b�~�7�>�-1F�j)�}^��:�^m��D�����r8�'�=��x�� �Ù���.�9�̺R�N�8��a1'q��
����[����RAA��k�����_��L��
f�bFJ�]�C}���� (V.C�@�YM��мI�B�4�����"����G>��2��v�*��
��.7��.E؀s�D�1Wc{vNG��������5I�=���{�<�}�-Zc;���J��卌�2��O\t�Ǻ۝�Y2�G���#e�|�L�p�&�Q�~a�����BA�R"����`�������~Zv� �q�A���nm��@��N�F���`���%<W��{#S6�M0E�h�YƟ�R��=��j|}-�h��:�%�6 8���N�|�|�H �oS��%�����B'᠐�"�˅/��bqPz���a9ϗ�!aȈ$�� (S��TA;Ǩt�P6�ѷtM4�A����Y��vs����Я_�=w�����6᪜vki�b��2��g�LӍ� �A8��
=U6�dw����
��1|Ro�P%,=%�hTUh����K��_O�@��#u@������+�Ŕ{!�4�f۫ӦOk�N�v����-�4�����-ȵ�C�8�ܶ���}q4��`���I	��'�TE�У��ƕ �#�ʴ X�߯nN��Ro���꺿��A�X����	����{5�^z�_Ժ '�Ĕ/B�MV��t�&��D�;i�Ǧ�Z:B��g�r~�)j��/�GN����ٱZ�~?�hl�|�k|�Y�Q�;R6�<�ǔ?)w�LFH�4ޣ�?��]Tͥ�6���ID���B��Ő~ԁ�q�Xg�q��3	�&�ޛ����]x�]��\�n`V�*��/4�TL�K��t�'�;�/:3��}��=;D�2E�%�8���!~�5�}�z�H�3#�G~O�6(�PU�o����z��&������Q��#�(V��'�4?�U�z�^�E�>��K�®�~�����Ւ�u?�`j@�Kd���W�{���5�F��Nh<��C�v/��E�p��E�(���b�1D��qγ��źR2����٢
�=����FdĤ�9��D�#�[]���k��i�&(w
"��'��̢����
.���,9�A�&���:]#�2qG�On4At��Xj���3�ĎS�*B�� "� o>i�,�gO^��N������a)�~S9(ڦ�P��
7s�ҡ�B�&�~!Jtʇ%��&�7W�b�As�:�Ŵ���������8�<ĩ�4��ȎF�;v^�Zg��;=eȌ�Pj��!����G��C� ?�\7?Ҳ��:�� z��鞊AN�׏Ɉ�P'*�����D�ť�U�F���|A��	x*+�I���y/#�n�ca��-$5�������k��ǻFnF�͕(}�+��rF�gYٓ�[h����5�7�{��EZ����W�%�j!�����x�jV8,������l��h�2���䦟��>� ��0x�̆{��>n��ޭ4�����V(�� ��B,�/z��4߲`�l�Y��l���sgb`�<A/6�E���3Dj*7TG�/��7!J�x;��HyFo���/��he��5' �2a>�nY���ACHlzn�\�{�ܫ��!&H��z	�(9+��-�ă��3<�
�_+�td�񋗽�f�<'݀WqY�[���B�TD?�S��_^S'@Z�.1���ډ������E�0W�t��������I�)(�A���>	d�����*Ѹ=�N%�Y���)_W)Ec#mN��W!iQd�c�^z�T����q�.��bT�y;Ә��=�dG��K�p'�`�J��xO2p5�gd�D�8�U��;�Sc�8B6�3�T^���"Hs�ZȔ�/�Z~��q(^KTo���;̭�cE;�0�>:Ւ����q:�4�68Z���BqV)Z�\�:I
���� qBu$<��pI�.|��G�u���״!2D�0z��3���g�S�'y��#��r��x��/�]�0G)���t`}�'��j�G[	Z�Ó������:(�ZG�~�����0����<��A5�M��2X;W%jX%q�靓���RqDA`f']o�D�"p�/q��9wHSit�w?�t���y�y\�Lь�r�5_���Eg:8ٛZ3ԥO����ufa���SE�O�P�����#J�,*��|Of�x�䄏�6HЬ"��ʽ2Y8���}?u���3%ך�����=O���;� ��q�n=�ϟͭ��H�0K�Co/b7��M����@�������wl�.��a�9�/~ɢ�[�GG��>Q�r��wyX��X-�-�M�P6<�Hg~�9�2댓���\l<��U���&�9�^���p�ǨϚn���P *B�q��7~+����O�Z�����5�r����,���T��'y"I��o���`Gd3��N#����W���ƳH�Jqy�A[0ߋY�����VU]�ȋ\k|��r��Lۯi-����g��P�]C|����W:7�u$�~�HG���?ݝ��Q�`�� ����U���,49���m~t?�u��r�f<�yö�Xp��%E	 I�_�y�g0N�y:S��WӤ�!)}�O-w�i��i�M�73qfc��<�K�m��%����",�]����lZ�����=I�l.Ŧ!��|�Y6��Ģ^�Kl�sT��=T.�����,A/M��ؓ\�QP�w}��Bİ�-J��Jg�	ʶ���X͖\���.��zZ��͵y��T�]�������ҕd���e=���w��w�.�l��'�#�Q�n�y
+n3Jbڈ���(z�c<�#׏MK*9��2`��_1�Ao�������	[�%��cɭ)UK=�ݒ����P��ߪ��<������8#�#<<v5pz�E7��z����I��"|�&Kf�!I~�E�wl���'èM6�~I��*  	�B�������޶�H]�ӛz1	}���ڞ\О^T�P8V'cb^�S�dR�R��~\�~8@2U�ƴ�szW)��W���mVD��w����M���U�����:�ƽI"�n�1Xzr�	b�G���%�4�s��r�x[����@?v�'���啯�&+����K�l��U0_��D]�k;9a���
���I1C2ݒ}���ì�)�\}� 7fm��d�I7q'Մ�al�eD�:�]U�Z�����E�����r��i͟�Շ޳w�#����D�RF]T�~79���x��_�
ȯ�?��a�Y���û�X75��n,7cE�
c.���(���Q�siG5`��t��н��udj���g%i��3��n
�H�Ȣ��������ܖ����|D���Y������1���{'�Qj�T+�e����l �#,�9v*�)�q��0���*6������S.C��g�A,�!5nb(�HDʈ"2�D�W��;+�whΊ%��H]�F��Y�D�S����ӿ��.(pk����P�N��M�iA���蝖$J�Y*_����'��!��d�����D�	�^�#�MU�x;!;�E�z��^~ȉ���F�\ŝ��+�k؃�@hOb��\\$U��'<��C���w�4�lj'RZ.��z�\�F݌�Ck(~�@2��p�)�#�zI�\~%S��5����uOYz-;�2��U���ȶ�� ����o�J_��Ε�-Ϯ�H�/�6T�!��%I��kl�	ʳ��h�K��G��zZ0�}��fE�( ��D���X}?�T�e���c����4����� ��c޻���?>E�@�����ى����I�q�:������on$y���Sh7
<eY��n��+Yn0�����o^��9�Ջ��q�/�HG��c�XX��}�_�.��q��bR55��yX�ԌԸG�I�·���TpQ�_�N2����vgua	���U��--h��2�{۠�Ap"���C�n��
ު�^3�ٿ���iXh���d������k`���$�2)?!0�����Dk-����#�≛ Du{!:8�?���&��ٳ�C�[����`���ŉD1��8�E
�T,�V���eR�O��M�C�B�0�s�c����������R�q%fP�m�U(�S �԰m�Lp���׋a`Re1 qp1�d:J�i���[�S�Wq��S{�P��]�����8�t�%`o��kV����!��h9!M�Y�WB���$����N��,5[�EAQS�S��&�u�c�l���^��/+;{����CUo�&����?���$�s�f��Ү�����C�S�+<���&&B��Iӭ���\�;)��������o\wcC�"���;x
w뵈���!�k��|h�!C}�gi��(��9��7!����؅%�oԛ�Ȁ+F��A�'��b���,�	�E#P��E�R{I�y̭��H�DN�{7�*��8��c����ݭkT����h���wp�C��� b&���+A����F�&?�`�����G<θ�<r[ܴ!i�lw2��'��f�3I��m���
o�Y����:�S�y�0~=�c>�*�]ݸߎ}D��rTI�G��@܄�.����j����AO���w���b/��,/ݫ_���X�3^���*�A�P��t��"���V�j� \��V���?�h��v��r�$��-�9��(�M�]�ƌ6?���; .t���Ʌ
�$����*���X��g���{��>^��z]W>_�.�euE������������Dl�֐/W}�j�vG�]Ɲ�Yl��/���<���l}`=]`xAU.�=�4��g�{��z�&@�Vk��C�%�[6����FZ��{ɩ�īl��{���x�r�G��!m6¿��:%[FN됝,H[=Ǔ
^S=��KWF0j�qml91�WW�&ybJ��|`��K��>_
1%�9�>n"bs2����S�_
�I�K2 4�E�<��O�4P>�	�8<�=#_~6z�(:�KQזUr��	�o�e&^��Q��j�ћS8^wbh��<Z�1�⊁��;�8�(֣΃��Z�,)��=��L�����3)B���jQ��W��k�K]�J!XY�.]D�9W�����"��/�\F(��цK�91�~�H��"���ŧc���(\�RO1X!m�s��}1��][\n�ǧjK��8�`������l7�����x��kY6�+^�չ�-Y`�Q��(|Ӌo-ɽ"X�� �os�� ��������hS��iT��g#��ל�p��?3�����d�=��u6��� i��L/��u/_�B�a��2n�X����P+	�X�ZN�r.��m[��%n�P!$�ޚi5�L����_��yy�a�E?i1�-�J:�Z/��F���j������u��4�0�ð]Y�����c|S�Z4K\E����*v=���3 �uOMҗ��V�i]T=�꧕��*��*�¹��0N�-e�d����:-���p�DZz�p�L:��X/Q8��{�\b�D�9�.���]
hjO�3Hٿ�����8�U�C�uY������:]��IT�u��&{s�c�P�,8B��a�U�M��݈\Uj�[��Vf�dLX� �S��72)&��N�� ��`� x���h3T
��ƹ�Q�>��T��`�ȏ�,����<�_�e{tDI!͜�� �9|TN=iR�=1���(�����#S��Kq�/L[��lW���R�z�Ш���c��C9�l��>�]4�Kx,MP`�k�|*�Yf5Ԃ��v���Տ��ncu|]�Z��R�N�d_�S�e�Ic�ј�S�E��70�����c�EM�8�)�[��Ъ�m/�a��IvJ�"%��y���4C��-�o�Jv�I#P�]�����k���
�R+&7�
(Ė�p�����@��j�� w�m��#R.�TJ�F���GW��C��g|�1�$t���%F �p&��
���¯�j�yQi��T����{��2���������"F��B+�Kn1E`����i��l�&oiY���}��5��N
g���__ d
�]C=TƤ�����{��:%M�T>P{�PM���֑�G�}&�_]Y2䇈.,���h�4��Ÿ��Ҁ��p����YYKIU�9��&I��Y�����TMzD�*���(E���T�=$J'��%:�Wc)��x���Tg��[t`.��=̛�W��P�њ 3N�����@Z�FX:�F���}�A�u�3��@�6�M6"%�O��6.��[��c-@C�����L=�6���4��c�ʟ�K=�������P�|�qܐH�������͂spJ�K҂�YԣO���w{� ��;����`y�����9��<S{k�U�F�HDd ��5ؼv߸C� ;��x0���A��m��"�&$����mbr����◾�Uܦ�EFt5���7d0�Խc_5���w�����E$6M1����x؁��wy�+D:,�at=6N���Rz�I�B06��pL��}U.�T$��8���K�U����|�%��e���o���Ə��+#�)�w(8�p��K������K魠�/ޮ�+��r���h�@�(�L�;0�KMX�*�E��Q�-L��u�OL-�&�_y5���9vfU˕3k:d2mi.��v�|�ܓ�L�h�,� ��ݑ�y֞Ȥ�Nb�K���;R����~z�J�z1=�tF8�X^�`�fqTN1�(Hk��{EP@WWڱ�1�o!wÔ��H|h�ck���_�8��iV���݄��ֶ� ��{�w�������XF�Wsr.�hR1���0�~�j�}�v.�v���	h6�r-3��Un��w�9�#E-wN��K����忊��������U¿�kv�,8stѭ&��Wy��\M�����>y�K�gssPte+����x���r9�D����&/w��g����!O�L�����r,��<(��t���  ��
��M��z�oH�Fn���Y��_�� N���5�%i�[��@]9L���©N�z;�.�ߴS
��/��Lf9>��!
+/�h�2;0j��������3l���>I�#U����{��D�a����]I��Fς�y���B�8jF��<�RS���[�e�!�{��[��TB��(Q�{��whJ�s���:b�
���Ώ����Cq��G4��?rhʅXr���`�eA�e��n��i!�R���]�{�V�eJW7,Y����JK�m����A�	�s9��$�y��a-	}�
�ƃ@F�["�:�##i<�e
�G�y�e��
��=��Ɉ)���i�|"��a�~�3f&è0Q�{�z+L׵a��0N|z�30�m��q���^pp0�ʃ{���)����t6duw�#��	n�6bN�:�Y�څ$������FR��[�����{�KJ�um�0�L;ڮ������H��#(hQ)��xrjd4�N���V]	�	1����s9��^l-BV����Du���RN��+x���;��=gb� "ۜT8wv*m�ң��^��b���/8ȶ�1T}^���m�K�w��Ý���A�UL�gN����G�N���b"����e��n���`�a�QŰ�L-b7`���;����ԖO�+� V/�[�on�u�L��T'D1J�*ýZV1>��<=z0�c?�r���qS���લR��P��X��VP�]���'G���b�=��{�e�jS�r�Sܭ��
����q�S�W �u1B�R[$�>d���uvZO�y"�4\���n�qG���2����}��z3-��Zx�,�z�ꭝ	L0k��R��}��(��!��{����9�x�0�Wܞ~u���罞k �$չN&��2kZ�?D��HϚӠJ�`L�X��������g >���^�ߝ	���?�`��LK�j�y���AݠKmm9wo\ӓr�`�Sϻ`��Z*\֮X82���|X��L�l�����f���l6�´�׉��bQShAjnÃ��8�f�,�%"�<PȮ�Sc�����{h�j�y���U��ٖ q�+�zg��#���9K�$Մ�����TB`�N�xٰ� � ,`C�AXW@��� �e���q�sT���^��+�Q��i��au�`�@�T?��G�t�p��.�s�����b�Y^��A�a���c*�W�a >������)N�����������<i/��5�с��H%�ߜ1��V�M�9>��a ���K�|;��G��[�� CuV7����y�	��Br� ~���E��������X�1n�ꊠ�IaqU��q�b��9�.�vTZ�q2��8��"G�Y՛�v+�<��n�8.8�0ݾ#�7�W0�Ma�>�����D�@zT��d6�(�o?��It��h��on;ʖ��>a}0�O�{��V�j�4�=(oS�B������@sP�b�r���R�U���8�i�wq1D�����צ����nZ�P���IF��>n��,��#�g�O<a��n�|�ML�rCv2��ȝ��[��X�R���EU�9���]m��i�[6R�$Q��Ʋ��9�Ylx�ghҀ�����H�=��hy�T��h�) R&��R�gw2F P�JH��M����p� ���,�[⫳'!�z�ClX������O!3*���K<()�j�H��Q��"զ�3���#��Ū)�R��8dC<�5�̻j1^�^0���2#
D@�8}�cҹ�+iʔ+��#�9�	� P蔰}�R�.R��e�z��!?!*f~��B��Meq�a���������֠m��^���4p�<�ZQ��?m��I�N��suf�1����NN��2�`��>��b�hĽ�F��r�s�l���m	|W/«bw��ܐ5�����7 q�r8������7��г�=��d�L������%"�)�6W��Oi��~��_�Lg=hNf��K��g�ֆ]��T��T����u�t��IP�+��	�D�H�-�+)&vk	��� B��^09���ѷK>�1����v�-�Պ������P��ə�=��w���b�� ��l�vS�z�&�Î�D,l���EP2O�nЃʼ�F.=�c���٨+S0���B�n�'�M��_7�縍UG璖�������!\�K���<R�Nn��}�g~#ߜ���+y�Dw�r�1����/�U�"�?p�cW�9��`���P�߇�ݞQ�^�єS���~%���|^����g�{x�)^�~܊Y�@�{��S6d[�g���tסm;��պ��]��E�Yn���-M@���R��Mc��NUۗuҪ����$�\Jx�A���0�L
�b��G���d�6�f��E���Ht%�4��Q�`M���d�������j�H�Vʓ	� �ĳ�K��\���*�N�	���� ��^�����l@��wB�q�;P#�5�r���x�S�%�^K�d<�P]�&8`_��M~q�}�>��D� ��!1���	g�����E��~a���3�ya��?�c���9����Ʀq�(�^�{pI���V6h�55O���2M7��^ �㫁��e5����5\o�-��.o�}��5�=��ų�_(����,
���}����[����8�N��uОC�ke� �y���HBy=�W�b��Y<�}"���/��
W�*ɏ�K?�tK�r�DcE��]��;�5�[���U���5�=ZV_i�.b^~ot�P_d��_+2$;���J�Q=V�%�VP��'��W��u�3)!�pk�8CM��Vw2��YC���f�������w�"9����d�Br�h��.�a>}��>IBt���i��S�6\.��k���d��JO��re�F��rr$�|��u�|� ����6k�`$�����w�>E���T���V�E���Q5j�>����>Z�Vq>h���� �YΊ��BV���8�-���y��6�%z���}�u��әYQ���R�:���	/���#���y��k��[X�e`^
t���i ��!70���C�˷���+�^ƭ�g2��
F+�NHK'Rk�~fߓ���a��G��dz?�Ȯ�ݕ���5z�T2������%�����0��"_�W3D8*�D%C�'�����oh��xŐ�t<J	�'o���I��P�ѧ1���8��!i<���h�[6+��0���}1��љ�v{�#ͻV���܀o�c���&��cIEg��sҝwS?E�+��� �5�3���\��%fFjU2D��x�,sm������UŐ����8�P�$� T�Mco�]N ��$+�ߔ���A��;Ѱ(B[l�"o��gC���'&�Bϭ!k�����{sAͥ3iD��P� �Et>w�ݛ;}�W��[7
�Yo7����5�1L��}��b�ǚ&���u<�]땛�'"��Z�܌�h���E�5o��)	��8���J��i[�ҺI��pJd�w0���O��-hv<�<vu~0"0������\c��q+vg7][�]\����]�*�O�N�|�D+���勸�
Yr|��HR��ӿ��ވM���LbP�Hn@�X�e����6�$��ap�U�:��܁���P'��`5/*��U����~.M�����T�wY���A1Y_�;�fո�M��x}��c�W
�sO�j�Vx �跮�Ԍ�:�"��Ç��i@af��):=} ���p�<M��\`>Z�hb?��<	�%��P��G���'���͛|���T��]ݻh4�_��j� �׾�T?��,2�mk��Θ�� ��71�'��Q@;,c��&�Z�n:[D:�%�"F�C�_�=�Et֩�ae�NU�#���&KA�{v��scw��ض[��`O��xaxdct�#�5�(�|v&� �A�շ�˱�z�T1nƋ��8�O�lU�JY�����".	7���>R�%�&Xg���sd�)�D�K���2	qv��~4ʴ�<�5���<c�v�B���i��}���Ŷ^�}x8Z���-��(��N6�
���N�_T��\c�?sǁ:���;5��66EFYt0��AR{���� [�pD%��t������3��8�>D�H�y�a�^>��T�-��#�Zi|g�Q�!vÍֈN�����<z?��CAFg�䶒=.%��f��%��~�{z�>�NT�Y�(Ju���r|^�Ʌ��w�<�S�+�p�1�p�o�L�zt������w(��>���A���>����m�ˈ��ǷW>ql|hÍ�z�n�r9������D�Ǝ�o���O�N{m�� �RE�*9�}F�VD���QA,���/$k�������í+���p���\ql�X��IOKD��X�i*=*a�!�bq6l�hZ�T]<Pl�W�?�R���q�l�Y�n���l�f,y������d��0�7�%�<�<U#a���8� �A�*�8�����b�*v=�Y?��ݝ���*����`��Z3�������"�����|O"�3��5ă#M$�Heg��H?wv�	*��jd��bXj ��(n�YS�`�~I3��Y:�3C��h�:�d2vW�@@�
<�a�Dz��8D�޶��8VѢ����+|ʣdng=��tֆ�1�N��zԎѴǝ�慠P[�O˾\�����0�T(3M-dV7���J͎���a�vd���]'_� ��֖��G�̴T���RR�5�]�%x��!�6�!��rHنyF���6cK�!�k�Օ�L�1���i�'�?������7I�4F���y�g`��;�{�����<�$�.A��B��'�2a D~�+mm���vT��v�
�ݯ�!��R�
c�'Ÿ^�@��._E'8��qS�q�1���
��,�WE��e&�K�X����W�1A����zVa[��֜x�#drJov�x%)�M��Q��7w>����	|ʹ/�a>�PӭȚd���]�(�cX���)��5�۩�F��>������PBB��<�����po�����8A���%HV�*�.i J` w��FqF��@<W��`^��9R��
%:��,���M�-V֚7����+]�{�8�� v`�<����CY�W|��w�ZB���ӑ#[ss{�2�9�z[��Uzȱ:1 ��׮��2 $��Ȭ6lU��n=PA�Chk�>،D���B�j�gvc��M��A���)�Z��{�*>ݐ�u�~M�h�q�� <����>�hV|͕����O��E�r�w(ҿ�H7m��c�e���NϾ������yx��~ U��qDO`Õ��U��f�ZX|��y�C@��L&7s.ޫꖱ��`�t��\������:p7����A����to����tD�"�"�`��U��~��c�4.H�|:�&�V�Kz-J������E�Ę�D�ݲ��={~��]�O5��3��`���>�p����t��_��u+X&��pw���0O�?+�Yx&��'݃��{����b� �>�wt��r��ᄈ�X�~���Q�Ҁ�f�2r�b�v��)y�`j.됿|�ie��R{;[��s�:�	Ah��T�H��!:W�H�����P&�N ��qﯱqqC\Sgn�Ȟ�D 	�>�|�=��9��E- �i�k��dc��'%uI��ƸK���(_@\EY���]��Q9�����{v>$2T�`aN"R�z�+@��,�6��W>��ʹ����Y�I�(���	�q�& :�C���%�gؓ5���
] ��&�_M�$;���	�/y��sBU�	w����0W�A��F�:۠	_��e�;l�[�����+���kp�nl��G�4����([�.��ˋE�H�&~a:���jƯ�`�"z�����.��@�M�[�!#���̆���Vm����N�U��X��_#�b^��tpSz�Ș�&*t�� ffO��cXCH��|�-�HN�mI��E櫽x�kj�M:9���N<��@��;���ѻ��-�}๎`\�&b��?�rB�����Ϡ>���w5��I�?i�!m�&�X����˱�"���[�Ǫ)}^�����#ݴ�Uy������@�
�~��{�g�V��T- �.r�^�]ρ�3r0�>�ٮCMfK�'��u����h�k�<����jj��l@Ȭ�-%V�Z �lO9�zn�3۹�X]�a 	m�'+��Hg��i�.��D?���)J�;ƯہT����d.��Q����Q���)�Gg^�uteϒ�)C�&���K�rn@��:��~?F|#��aKX�*^�[���ʲ�Ud}�kט%�L�RQ%9|Ӌ���T����"6���56ȖR~Т̜�!��-���-8�����醺��$91����X�8�j'XN��ڃݿ1쇼V�&�Q+>�f������'� RИZ��q���Լq0�=�.fi�� �ɚ�c=��6-�r̴q �:T�G�����x䣡�@,=0��ͥ�E�s�(e�s*m�7N����Cw�a�@$�_������bl(Z`z�e��z|�1��LPj�y�k�X��}HC�&���[�y�a��G��\��Ś�M�k�k�M2;�nov��Xo��I(d��'�:��D�(�I����~H9@X��V���.�p��W7	ԗ�^F|K�#�>�֑�t�M���u*�HgJD;�C8'2�Ϙ ��ZRW�l��#�6��躽>�P�Rz����%��6:s*&jO�N4�廃iq񾘅�N\��# ��v�7<|����M0�NR���W�����('��������暈 ������d�	ץ�����!�����Y����K�&������9uc�ը~�[�υCk��>�&�M@%TΥ?π�(�1L�e���Ig�2$����}�ӫq嗻�ڊ�UHok<'�-�UcT�����{��Ə�Ced�fH��>���{
���*�:���6���t7�FS�����-�tޘUfo��������@^�7ql�*����Y��+� �S�@�=`Jl;�~V}_��Ք6O�t&�ה1c�JaȏR�	t�3��`,�ֈVz�]����1e�q��N�u�8F��� �@\�����`/Nl�)�*���m��"�����BS�&��������������	�	3�d툌MOI�<����d-<(�:��T�iﱾ�'m���r���ЙsF7�Y��@NMI�"v��ێ��]�'?��4�<��̋>�
\'�ˤi6�i(�{1�lU�e?7�3x��l'�`ӎb����4�{����	Z�T�U���t��e��A/��;,W�=�<��X�K��)y��T���˵T[G��Uw-�\#��������{��q���0?φ?������s4��c'^�L,�Q��3x# �w
ה+e�؉��د��F�tFY(1�%���;7(&��x�;���.Yi-gu��U| ��h����b�	�W_�!��m�l���it+�Hr����o�A�����7B���h �]�r��#���z=�3������Ȱ)�t�B���s�G�}8gfآv�-��2�op��!a��`q�)M�~�9����.E��l�(ܦ$?��CE$�R���[�!�j�ruӘ�6��@�K�D���.<8��ap�rc-�By�Rm���P4�cʈ�Er\kT�~������ӵ�x���X�H-�)r�
D�ԧ�s�	w����i�<&-C�@�D�J/%{ k�ZI�zX�����ӊ�@��s�������5߼s�#9�:o��T�wL�5A��E�#^�����2A�DX���wvͿ%C?��(�myAd2�o����lB��=4~����:
�w������i�MV)m��'e!�z�\�knbM��Rsڼ:XK�;��7���J/W�("��1�QL�gtT�a��]�y��"�e�x9��*���P�AV=`� [f��.��0K�7E������d
����j�nP<v�r��	9�F_�r��YHw�����Z~0	�l��rz�`�^��8�Q���P^D_nG�h#N������0fqO�O�mu��)\/ ���IBW�t�c{�!q�{k��{\䥴�n ?�7��:��8��>�TN��'�_Y�/B�z�V��i��&���f�;	W���U�@�;�H�l�o�M	L�0r��Hg�Lޯtg_��j�`�C��+,"�5���}'���,8��	�M[���>,&q��~����ς������;t�i���YU�Yk`�Q����
YPh'�^�7K!���~�+0�j��) C��ɻ7�j���b�>�澌�[�!�I_&}@l"	����hĘ���t$�i3_��U�$�&�W�_��~�eĒl�P�?�M��#פ�5���W��x�#\�#)�	��A��H�8��xyl
���,u�z�	����4{�4/<5��&�v��ɱ	m[�癅*�9�Xhg^�D�g-�'�2Q+K���@�հ�B)Ow�La>�-R��k���N��T��Q�'�cL.z��������Z~�V��,M�~�".E�d�:?]�GO.L��(" *cA���m��{Ot����g�����mHO��E���V���C��@�5`%9�+��c�B�5h����n�\+ !���_G�]�I���Iʿ:T���Y������Ōi��x�pɋ��l�m�]�Z�Y�a���s�@b��
�M�ɯ]
Tb��5���N����W��^SM�z���uV��
�J��X�}Ygj����;���D�M��x�Z�dS�,�ҷ�g�B5����J�P�=�l>q�]�yӼN����cw0A�
xM^X�j�3u��y(���:ٜGfu'����Q�)f>��𦳀�/:5�$��J��[,%c���0(��Ӵ�r"tM �u:�N\&�����^�T:�E�e���L�ohs<$��D�����L>�-k��s��C�2�6�*��Jd��vKXH�0%oD��J-��`�2�H���	 �3� K����d|�F�$9��c�ß��-�{�:������J�����Ӱ֓�f��k
��oP�5��3,�|���J��,k/��aB�ZJ�?'n���V�[�&a������Ҁ���}xZ����X*P�
Sg��g<�@��������5�_MM�����Ae:b����N)UZ0DP9RLA_wW�<"�}2]�:�؄������L��tgj�z�s�h��~�d��c��Z[����ȝ��ch���2��>�0�V9,h-!U�D��yF�kr�l�N�@���^( W��*ag����4�i�Q����q�Y�Yy�>"c��2�S�E���^#!S�m�{�*\������0���4/�9@�a�k#�� 
���~�qw,��!s��cQ���UӀ[�1#�Z !ݥ�I�#KIc���[߯V�x�-~<�����W��A��gu�����C@
�3�*��������M�g����z]�G���P�� ��t�� 
i�c�t�}_b��6�b�O��ŝ�9Z泾!�6��oT��&bp��	[�H�Mt��g`��5dg�6e��O���3Y%��<C�E8x�ULg!:���*��5Zef�#�0/�&]$���O@�ҵk�X��	T�E����T��ːt*V#Ěh��!|�)��h�tcG�R����wHl��)a�Ie��%����q<;;;�D���������D�"�V��)P��:a*ʫ����J�Q���g*��m0a�U؋+���A�U;u4�h�5Ӆ�%��w���9{*[HP�n����%�^6�%����QXϋ��L�c�v7YuĻ��Y����	$�*��n��V7A��^�V�Q*�j�µl.�A��^!��"��`����J�܄��V����qv"��dy�����^�e��k��-�;��<_*z=*��h-���u���d�t� �j)G����P����;���X�@rj�������pO���(/�?fj�!��ПQ�0�.� �( �\V�%P���V �#D�D��> ��X����D�E�}��dQ�(;yA�%��f0�s�0�e����Kj���C�VyM<� 0Qܭ���J��GE�Be�~I:'7�\U%o�*�P��	��˞��us�DE ���M���/֩���W�ދ�	txC��2�i���G��O��Un�#��+�e�u�LG�K}Gg�@Gi_�� �h�7�#��/w���\�}���I|�^=:֯�'w\� ry#�/�_B��)��g˘��3[ʯ.n%w���x�{r��Q$�����Z!�aH�W��&4�t�MU68p�V��4$��oަw��ݲC�3(bڕ*�D��z���	��h��a�cg>e#�e�h ������ W��b�EZ������O��/�[\ͱ별��Gm"���?�{`����(Wd׹~�6�R�Õ���Fs�rx�.*B�!@"<�gR{�/|2y.W?��8�E���#�vc%"���<�h���x����#���BE����hx	�o4o��J�GR�r�ESgG`7��X����G�9@f����"P\D8&��p�� �P�j����[���^=��̭���ƭb�o�������X�U�D�1��?E�XNW{3�j�f� �@_~�|��CNK'T2k\`���娸��T��j�:�h�F[.9�?n\+ ��I�P�X	}�qs�w��)�A�`L��|���lit��sm,d]�Y%�X3!m���[̙�:��e�Њ���h>*�����FZ_�ݳx�O�+a�%3s-���b>��ELCL/P��ɡ+�m�B�g�vU=�\��	��5�N��
�LB���1�a� �R��d�%��|d�VGP�l��(�uoj�-4>4/���-]��[�0��������SK�B=����w�I��G��(���"l����ovY�/����n
ֵ�p���h�X�|���c]̢���Y'ni�ծ���#[��T8�t7�NV^l
r-��_�k�ο�����vG���vG�1R���2��f�R9ᤣ{KK���5Hh4�?���,/��qō�h�͘^���DGqh�����D[�"��'�EaȒޅ�(��4X��B�G+:p^���=����i_B�~P�%��a�x}r;b�NGT�jAWrɣ�<�I3�s�� ���)�����*a�e[}��]8н�x�3v&"���Dӄ��8�&
�B���.0|~q�5�D��+|��v��w%�L+���|�i2e��v��%6TD������kj����[��u�i�9_S�B�Qۃ}��� J�DN4(��C�ja��p�Ru:t^?���ѻ��u��;�{آdA ���� ��6��b�Zp�P�H�[4��,nF��.p�=hl�	r�QR=��t#O��rd�	r+�6�Is�������krE	�ϛ0B�K����i�T&���	#�糫��1���g��@�)9�P�I��#"ȢW�uN�I��IG_"�
e���G��?(֡˖�Y9?\�W�� 7������ xߍ��}܁���M\i�OT���x�w�Ǟ��xn�(���Rj�r�0k���	����n��~�g�T���l�:�i�{L�V��[���N?�Ob�E�{��?&���	��Ҟ1p�rS�C���k��GE�FN��
���tb�	�~�"+\�{�����ڨX`�A������f�;j��X3���|mY�ѣ����u@Y��MH��_"�d�O��z�=����T�硼����;�Fj/��߇֞�"^k���_��u	봴��\;�����JNE��G�E����O�M�����"iq.����#�zu�9z5�~��mUGA���T�@�a-�u�
�`�{�Q�W���u?7	\�o Յ؈��o���b�[�&?�v�������k����G�B8�c�26ޒ`��}�"8�n�rI�c�6�2x�|챴Mh���HC�������h��k]�����J�Z�1��h�c:�ra\Y"�J+\ⓛhE-E��_c"u,+]�>H�nm��ڥk���O7�#�-(�4�Ԩ4�E�d#	:l�װ���R&�5�]'��{*�-���_�Sp����zc�a%)z���S���,��D.&�Z��	��R��*Tx���bf"c��Ie��86�'��� ���'t�
g@W��%����%1 ���b�P������st6�r��������M�<��M�k���x�8Ь�:�Cè�|�Xp��<��'�<��x��d���ȣ[ &�i_V���ȣ� ���c�rBeߠ���7�.B1Cn�u��t��yVR��'g
�hڭOF<$۶��;P9Zc&O+~"x���PMU��NZ߷��C�8h]��ݩ��+�j��)bL��ZI	�O�iA0�n1����,R�(J��js�l���XR��]ܘu��U'�B���M����	�tiPeU$��"6�M���c$?]�ÔY�[JUIڤD��iM%�{��6�0vϝ�//#>/)�s�~A[S����ɵ�j�Y���lT�S��?�H�1xt$�3�g2m������(.]�>Un��F-��~�#-�>M?WAO�e�^�e��x����HN>���=����!��(f��M��
���}e��-k�Lh?.�G��y�󏪿_n���|�_L|���Ǒ�'����V�P������1�;'ÝA`�iO����u�^kӖ�u�8��C��.�X��D���r�4�b�[ɘ,��r���s[�	c �w��gq������a�)o�Շi@�M#���R�%u@���c�����'d�:<����1I��W[7���$\n�g���F��~R~����H�����S+y����s�>%��;aE8�5Y �Z��:�G� ����j`�j����U	+�,�1��V���x}�$X��b|&�3��9u1r�4M�G={Ԏ��2���z��޶�Ogm���B����eq��d�	�R�pJ��Q^��AM��l]�-�1�Qe�N�coN��O���.���0~ɮ��?�T�0ٷ]��Z��)Х������p^HW	����h/�A0�0 �C�4d� ��7+�=�.t׸�=
����=���4(�6���{���n@�����-=;51�wj�9�S3�%�0�s�c��@1<)���;9����U���r]�7�]P[���Ug�?*���7h%9#��]������nW�= <,���M���5���A5贤��Ċs�������C�Ձ��u0�\F��D���<5	V@>�(�|�c�	�j���I)���?Db[��+c����@�4�}�(��2�_���2I�����jS*�?Ф�H|X��D�Z�,�$$��2M`���p��ڳ@��U\�����ճ�&0 'd��MP�9�R�Ȋ�J�)�;xh�~C���p�5�����to�Wo�WI���|���Ć*S�P� >|nt�O����B��r�� �\;w^NN�L���Cz7�_@n�|���7�`��"��[ؑ�O��v�~����+���+02kh�wR15�]y��,qa�d���O:~����h8�3�=�0����fN��?����i���願�&~lk�#��y�")?C[t����v-�H�����B�e~��NB[f�T��X��Q���Wđ���d����Rpɐ�p���A����Gz�b����(>�Ǔ�A�����};�ӎ5J�K��-\�C�	^�
D�;V�-{�0��]+����6]x��N$&';�nJa% n��.���prh�^Z5��S��������L*vﭷ��'��O���t/�`}fM�����jʚ�8�<=-i�V�@"vT���
���&�=tC�4����&�P5� '�w�(��$ΐ����C��~�\����D!�W�s�Ou���4i��AA8�iD$0�1��(IiGs���ra7�1�ױ��/c�=M;.O,5��a�>,��� DW8���T]��4�^	�ɮb���)�~��i��b�(D��O!�bn@�&������m.������8t������#y���9M��qgs,ob�^�$4�L�g|���#�q�5� F�=q�o�>Ίx`>�2f��^��'1pFI��*.���6���}m+[M�b��"W�E����	8���݀�����h���O�C
 ��.�������~��^�W9z�~�reY/O�x�;:�;�8�[/��&���l�р�y���=�����f�Q�l� Sc������{;Ԉ�ݺAq<̱�L]��]�U��j�p-*���Zw���)a�e	��κҌ	W�
��a1���oKK�خ>;��1��_^��u������Zt-�C�gw0k�xI}go��56o^T�Cܷ8 �7������;=��W����=L�� 1Z����Wo�4Uk�q������3\3��6�)�oV�{r!O��Ӌd�!�cJ�j|���=\�e� ��G�P�^aR�$·T�eR���،�8��)<q�͒:��-�J���1��%�п��k���}�6\�O��MC������H�	خ����68 ����X���XJ�/4ې�r���M~wIu�=sΡ>W�:��m<��l�u{U�bvf�94�Z�Z�r�+��tc���?3���+>=�)Oo&o���j��j*��Юl���Ѓ��];ÔX�`����̏���]P�ѓ����+�Ȕդ����Ny�4��HD��⯼���Z��+�w_�;��%tg�"�`(ް��<5%g�Kmu���MsZvOq��)�;h7��}t�#�%��6Û����Sv`O����� �T���Z��"�?Q�R�����:�����m�<�����v�f����nK���+K"n ��B剰xF��<� "Mv�+x� J��ǥ�;����@��^$�]A������qb�8� 򃍫y5�<�c��U�d�����N<��P[Z���{��"�qy�9i��a���E��,�[��i<.Y�w|�˄C�M1���݌zgz���F`�b9��?Pl�ezՐ��P����DY�F�����B�#����o��m�d5�5����\"��m��A����2� ���u�@<͠�{�"a�V��a�?���+2��k���8_�_I���u�HĚ�|�BQE�Qd�*�0tB���1��Q^�����(��Ң��w�H�pa�WI�W����\w��$��Z�5<l�M�A��j�-
��f}_'-����<^)=;e�e�Ʉ��>daJ4XXnY��rM�-Y
�u��B�ޖ�58Lw�npT�u���ᝄ�(�c�Ex̑�Qlvo�z�D@��Q��<�<٘�OQ:=���="��3#�G�"�]r[��}���lU(��fy��y�6PT�d"��<dX �KB\�����Ȍ���ZY_L��K7�ʩ�\�lC����)t�ϰԲ��'�����b]�|6���k�akJ�k�D���ED�5���ubw��2���@�KDMj����|`h�`\�"a�"eBk%��ͧ�-5t]aw����i��J�'�&u����ҭ��׆�D���%N�\����!0?��r�h��?Z�@_�ʯOi���=�UMYK��r�3v���)~]�$��L����\�9�
q�M���K�bv4)�x�lt6�f�ƀ�zǳ���\�� ��ԇ4�l�6t��,>Q�e{�y\7F����������ο�c�MA��	W�C� #��~�� ��o@t��bO�s��h�9�g�\/�9Jԯ�f\��;M�,�x�h�{�J� u�/�\��UՂtl�.�Zsf@�$p�ɧ�N�1w����� �A����_p�7�'���ǵF��8�>���.���DD��\��/x̐S;����"U�*ڭ��0��O��Ѻ�lY��J֌x��H��+�Z����jO��l��-��(ڻ�A7����Þ��m��A�uȻ?e���~�*����@�<�+?� }r���D�KQ�h�.)��T�;�AwG�"lL���	��Ʋ��v>����n�ˇ��ԅwt�?PTH[��3�x
�����s�5u���#iA*u6Ű�"Z6�7M
i��?O�
iӁ'2��g�5��p�	W�#�f ��!���G�L�f������î0�BLX�w?)��\�YW#E�W��EqJH�x�<��P��dW�^�_�o}j���V"���6X%'t��P��Widw���Tb6(bY�NT���] �U~���MDkX3Ȟ�$\J��3�Ð�C@��e^\�'��|h?�l���Z?����z�R{�x&�k������d����W����"G5p��艖����8��<y��k����-�%�6s$��*rjvD��v�j
}�)3��R�/l9dӖ�g�RsR�J���C�I���a�p�ƼASd�-�#�AR��-XSR����r�}���_'c2]9��K:��S'�yx���{/�f6W���X`i��Z��5@����;�*���|Q1Jݝؚ?�D���ݍ��g���h�*]f�{~U�V�Z�d�Z�(7�ZL��&�1����4�)�
B�35��=_Ez�e���v��B�a!{B�AbW�!�A��R���d�}�)@Z�����2���qMʁ'�[,�g����A2y=��k�d�o�@^(N�7;�%©w]��(��	��D*��^+��*մ-��(ؑuu5�x0+�T�gy>bx	X'@6�lr��*���5�{joNv`\�����������ˊG�x=4j�_�'$��׾��+Ky��h�]-�\FVf�|��!3�t�~�w!چ���LڀGr�f�)<cd��L�@�� `M�-M]q��FBK����؉�.�t�6��S��ṑ����	I��
J�����4C�9��)�-ʔ���'h�V*B����|BM!A�hm�)��Fr�upK�%��1ov%�|�IT1�T��z�V�ƟlUoe]Q/�� D��T��)&7�y�"�۫�2ֶ�\]pz��������� �r�*���TQ0?��j��_��%:/^c$%=�௯�����X��y��U�C�;��ݒ4�N��I8���|�ޟ�L:�UΔ�)�ԗ��� >��}��xE�) >a۷s^�Fv�[ˍ�e� ���$w�N����v�wˊ��BR����3#X!Zܽ���qA?nB��6g|�(��e7��&���cV�Vp�����9��27���޻~0�r�$�C7Ө�hk,w�#Ik�%UGWB�3s���s�u"L�a2��(.��?�j�����I�@�+�[��~�����Ĭ��Xj��|��h�z��֠��� ���QE�!B��Y�Rv�����Zx>A�-��}Ô���ℬ&}q�s�ָY�1�5?��g�%�	�9Y��T��1��jz3��l-O��57�f}p�Ov��o4���M!|�vC��i|��.��i��kyXxK������k�3x�������P�'uxI��&G��B�ؾ0W6���(;5Q*,��=�,s�-�e�OiaW!�N=9��s(�Fy��f0��; ����V7F�4�ۊ!t�R�2��{��4v���_�~͎HKx쒑�b�����>��
�j���#��Y胵�&��x�}�!��T����Gj�Ɵ]�O���絮a�S�<�>�CJ� �;�}z���� ��R�fJ����qewL�.���?i�a�9Z`<�G�~�� .��J6IpL�4֎Rn~��� �n<�È�^��;��gݠ�o7>8��c��;���u��fB�7ܲc����\���(��M�4������W�A��+���%����0�s䉅�+�胆7:�']v�;�� fW]o�&ı�M9$B�⵼�����������f<Y���f�[̠�Dd�>:+RDK�R���r���!��J�ThM����Ý����M��P�7��>���3&n�
i���H½b W�J-�}y��W��ǟ���vˡ����ZL.��@K�n3��l�@^��339	��3"�Li0��ͻ4>�:bJK�!D���#E��J";(�l[l�Rh%�sWS���<e�ZrX�B��3�AV�X�@�ֳ7����h��3�op����BBD�X�っ
�x�^���p}Z���9�����(iP�6S3���*��%���;hGr4BQ�%g�򢂨�R�G,l(���
;�_癩�3���g2�9��f�ÄV��G�\?1�N�e�VH��l,پZ�� =w̳0�x�	9��B=�ߋ���e�F��ۘ�A��
�,�I4��b@�J�y(���vٓk>+)��]�WU4�
�,���.%$�w�#&V��-���Pٹs�w߲ؔH�C�q���a�TGo����G�G3?�����4M�q�_���?^��;�J���:*��LPUHwo��t���YU;�RqB����#I��SY�2��UŘ�*���w��J�~n�4��NŽ��aih4����i-wq1�i���@����-��P��_è�)f$���E�	2�-�wU�Ƥ#�t��ir�e1�xa��D֞&�r-��Ė�/��'��{��5Wgt'�lԳ��LxB�:`��*$���,!��=��kv�q[��J����:��ВA��r�S�M�JKZ#��3�55�����ֲ��q�1�%60aT bQ�ј���W�Ev�M۞U�pX-�=�@�Z7C"���T
��	8U��s��lE��� M�=��p���mj��pP	z�a.U�5�j�$N��*�*����1�Ғ[@�1�0S)q0�;��w��qK��c�g�U��Tw�#*�/F
�j0��^i�jit��?2�_(M���;�_��+��	�X�2I��J�%?��~�q�Ϡ���=�J�4�ήt�W<�����R�CZ�f ي���31h����l�ЫL���޹�\<��'��wԎg|�{
����ILphI�e��=�PvU�"�?�&�-���q��/�ar(�b=�0�� މ壷��ɩ�p�dDn�+��q���6�R�F��v^�*��NV��ߦ��0�^�U�G���e�Ww�Tc��P�ؤ��"� Ql�k�T���be��FՔ$~ߖ���v�s(�b�ҊR�8��ǯ;�|�V��?��)܃`��W]�'�K7�t�UŐ��b���)YAm�a|��CgQ��}c����d�6#ū�a^�{:S-��4�f�/N�h�uD����g��p�=k;�D&�Ս|ۢg�2�:��Z�"j�S�T��pI:6��	�V+P��^��j=��D�M7r��@p2��>S�M2b���¢�?�߿��j�e"��?�L]�48��'�r�b���ks �d�����{ؖ�D�	�b�{����V2�"��v�����u����!�l$�Kֱ�(/t�>� �̧x�.ܩ;�V��̔K�"LIRd���D&�������h�D�z�n��5��s�a,����wP��!��YTF�tY8�
�h�O��������XG�%�չ]4�ڄ�h�I�s�E2�����:�����}Se=���n�7��l ���v-?�Wߍ�·�����l6��6
�2 �o8�;�C���'=܀TQi�RJ ��h��<	�+�鍲���]�:���ৎ��!
�;���r���F7%��ߝ)�����+�Mx�������{������������l�@f���+--�J��-�}i������ni^�#X�Ǳ�D�\��p�_vF��e:���{
y�nN�� B;l.��9B��(�ʨ,�Cgv���E��Y�⏘ ��~��"t����6t��%/�_>��*R������`��㙬�M]�K��<i��,1�o�����#Q�ahq��{�C��c��B9��?�#�y!�)e4�|���s�xS[�#��`�Z�1���T�R�F�+��l��᷶Af��6�\���6�~"�wU)�:�#an[V�JD�����ڂK1�6���3p��1�$U�b�wgM��G�a!歂�qȥ9{�� ���f�:]��m�����~a�w�b"�7m���ܻ��1,d�ʟojh=>�^C�+���t��gS�Y���u4�v��L���e�$Rv��⧕���n�@�Dl^��-#���&���`�>_@@ӊ�����q��ό�)����?���Ksٮ�$��.�n`�B��)<���J�t�1.1'��W���&bk�ԯ�����~�;8M{��#KWg�%d��_>nse)�6/ "C�u˶�д����,t�����0UYG�;�>̞�)P�]��ga�����D������d�t]O���6���SN2��D�O^_dl�i�D�BԬ��\��tH~�䆁*�" ��ܬ�l�	DΞ�0���@�L��E�2w~�)�o"f__��B��!��֯z;��VN���o���vqB*�b">m	��|��Hd��b�(�� �3@'ѓ�ɫj�ίjZ�����* ���/-̿�m�U��_U���m�	� M6�x%@x��,V+�[c9.m�6�<�[�u���C�[�
���븾Vxw[N=K�6%��5w�/�N�������8�Z9��,_M�hJ����[8~���K�7�C�VѾ����j���R�"�v�)���"nqd�C���h�a����T׺�}{\����7�\4Й��q�l&u��D2fU�<��c�?]��;��L)�p�k������6�Њt���3kvQ�/�G�G�{���S�S\��M�	��}ة4<&	d}4@NKز~��� $��}�i8�򊙲/�ż�s�8�)�����Ej��=�>:���{9����cx��Œ�A�Y�w�����"mq�r�fhe=�>�qh���`!�����nN��w�IZt��e��|���v<��n-?�M���[��y:7�8)^L��)Ь�	I2����U=ET��Fd���?��5Y��%�W����m��C�]ߪ-Q㘾���d5���ʒY"dc?����{��y��8<OV���?�������}͞�5��;B-�_Hd8>�W�gs�3��������^X��ɉ1�zU[$�Tػ��A���������FB�N���*nș88�\��Eړ:�lVPY����E?l�lZnZ:�
Ʀ�B����h ���T�Y�b���Ε����0'ـR�3BT,{#�	�(!�Tѫ���=-��~b���.*P������.�e��E@	�E��r��<�G��e��o��m�p��̍hTw�88����/�$=B��t���C4�ȑ�	���Θ4@�<f��Z)�����*Ƨ�&��_��15m��A��J"�M���;$���Y�i �2-�4�}⍒mK�b�t�������Z2�R� `��+d�Z�d��H�6p'�?����1WD�AA	w�5|3�*"j&�{�ZV9�n�{,S�A�?��n�D#�x�1�R٭�ӡ?�7�)�ͽo2W����<��(�`�v��dq"	JQ,X�b��0{ަBϺ����.~�5t�qm��F��%;Wz���D�ICfV�·��3J��[�F'b54k���#Rl�f��
 b5�f�o����.�!�P �ͣ���@��3���i6l��ЩP2;Ç	|�& ������_3��k5j&����"��hO/�O~�կ�����X�;N�QФ q}����8P����W̷C��ʸ�BpR)�Ij���V�}�7	R��vV�f�Rf���R�o{��qcO�vP9&�^MW�)-9U�P!$z<���>�"`�mK�h`9J�_*��k�j��.�/��Q	CO��'�*Ӎx���5�I�7r��p4	��85�<�W��t���P?N���2�� +�vm�`�ͷ��Le'=y�퀵�;`hES�Y��Z��Ԯ��U�&2�~����MW��e���Y3�,���������T[�p;.�C!���~Ś�b�U�BjW�*�L� ?'nw������%<�l58Hܾe�Z|�>�XY�5��I�&�z_Bd��ޭ��43H��TOc���ל�� ^�x�u�͞6䆎h���%D6
{''���TW��&؁��69H���4�Q�&��a9~����f��Ω̌h��2wly�+#l��^�VbZHJ��k�m��D���'�hI˃���;q��u���ms�,Y�����ʠ|�1r�'F+5i�T�����
����]v�f���(H5��ɏ��n��!����&�4F�V�$�2��U�*�i���ü$��_��Nd@��%�����1J�	Q�PE����0��|�ݯ磅W�~1qEb5��Tg��:? t#�Ӥ-
$]!25��N�%F�*���M>n*�e�P�e�YYW,�)E�0z��Y7 ~I��T��)s��[�c�A��'U7�1��k���K=#=��}����׵���Ǖ��|���w��*)��ob�#����_��5+����M�S�I�Wՠ�v�q��h0�r���'O��ś�����dOJM��р�r'N�}��%���D��*��ש��鰶����<C_��U����g�mB$̇H���r�Z��J���:b8����^�Ģ?��{�V�&���IT8rFQ�J_�m�P�И�i�ڥNi� Wi�oR@x�nCw`��?�7`K�"�oǺ��`D���V�zA���_��xe��̬�Y-��.�Y�49�Ԫ+t/G���u��kQ���p�EFf���
v:#�+�7(?(vQ�"�������b�q*å�_�1l����л�, x�͹���3�ę6rm����QN������7��G�!�hbX���J�|�����5�uV�5�^gm�|�3E�!Ѧ<u�rY����(=0����ݬ�ݠM�4$d�O;�6��J�G�K�[�	c"p%Q�"ON@A�I���H��Lc�x��1K��g�S��ӄ�t���_R���=,e"#�$=^f��AN,��ӻL�bE��8��_��l��AT��]����7h���rTaQ������"rfNC��y�K\M��_��'�:+K�a�F��,P���/9a!Ă�J1��;����n !���zQo�gr�g�β��_ ����h�e��	�BB�A�˂������ѬP�w^7@���2����~-��)���Ah��Z�mtVî��;�Q�3������)Yr�<y�aTE$ ��]�&�z(!IƏmV�ȠHb3�-D(��	%�F�xM�r��wΣ��ɜP1��p�	�S��Uye��� $wrK$�F"G�/wv�qtɄ#@Ս��Ub����p#�E�  �Iy�d��[��#��p-':LX�C,1��lm^�YQ32���\r����Qm>���Fd\���;��O�pD[�i�U#��9��Y�k5.8�����g8R�CZ��S@&�U�M4�*2��r1o�U;����F���Z�_Ɯt��^�wnDv���R�~����r���O��OҒ�����ƒ�AI�I��8��¦)8�2�A# ��1�q��B�Q[����) �N�7�FW����AL���[�F��/vΕ�|���0I8�`�ė�.�P_ƚW���ykK,��ތ+��iO�����g׋���#T ��_l�1��+�\ݑ�9���SU�� ���YxL#�ϐ9�	�1owB�"�s�@��=dF.
}\ r{���f�Z�S������ �\E�����u��Z �p����Xg*�b�a�V&Mבџ�TE�kfs���pN����`������zS��J4F�axή�Bz��4���|��O�ȉ��Ҕ�2��R��3��gV�+����"�ͯ2'vB(+�V��[�t1am�؍d��-/�_sK�TKπ�� ���j��TNp�"�^����dG�eZ����X��γ��vP�ƿ].L�����Ij���qV�Q��?�����#�zIlt�)p��Q��,������!6�q7�f��"۩�]�+���Éu�,/�?Ë� ��ظ�YF�5��B?av�[�ÍH��r&�=_�tˉ-In�^�PSÕd:812�?�?���T��\�z"���dt0i��5L�p�N[a|���cX>�X�=]2�%>O�lV<K+&�nr�|,�Np�mvb��.?��͞�fF�:���KAyҼh���V��D�\җYKUi�0�[�»�ڗ&i�T�~v�4Β����jf�H/j�U�V^�۸����F�����V��g�Z'�����k�9���=ˉV�A��> y��ݤ�������8��UBbՔ��*�G��W!R�/�pn��bvg.��4��PA�$�f����h�����:li�`��C�W��L�̬��s��C;�@K%e�x��g�(�|����$���u��M���G�.�9���JhN����C�&f�ˋv�n���V��ឹY�����ٶ+���C��@ۛ$�r�5��b%�0�s*���c�Ǆ,U�h4��ܦ��Ĭ1]&��>�Wp!�{1�:�7�PI7Y�R׿<�G��W�z}U�~�+ ��$J���+���>�(/kd⶞�m�C$(��1��o�a�iu��ː�!bZ��},��᧪���[�9ZX��q���#�f[�-Te���;���f�5�޽!��d����fj���C=�3&�V!�B�K���A����p��I��_�_������Vk�#�y�'
��a3$N	󱂗�^pn��X�M>�Zތb
�yp�v�Q��-*W�4��K���� Q����d����Q e-Hy�a^���TP�;�������8�c����鳩�:����CmQ=g,�h��P����K��)��������e}~z��F"���Y�����H��DZh��=��?m����[�̲i�n]e�z7�6BXR1��\h("�=��>z�*�-IѝX�id�F�]9*o#2:F���y�tIz�2�	�R�����疬A �I��f��l�X-Ha�iR����w��X��!_}]QPCzu���^
fM�Q��;:'e�%�>}s^��uwq5�ő?��#����F~~M[Oc=��\,���$:k�������1�zS>j�C֊���eP:o�;�]H����k���I*t����`�����xՓ�'��wq�kʠ߶�6:���W��\��ڽj%��}��x�K)��t�r 6�j��К�d�^B]�C	;��̜�݃�>ܮ2�n2.�4��P�aWf=�a�B�WZ��C��L�T�F9+e���,�B����j����FbV�k#K�39��W�$p�	�S݈_^��Ah\���۵Q�|���h{qŬH�ƨ���ػi,���[�v�w��z�z���̎�s�Ab�k�$8�-+�O�w_�=)�RZ��YF_Jmw��)�@�dW�� h�]`�����	9_+����.h<��2�<b���y��!�E��5A���Շ� "����i1�.7�ee3���v#�BIX$V���T�8���sӔF2�����l�f���ǧۀɳ�j����칕��,���B9�䨑X�� ����p_�Z5 %�'��-��08#�r?�ڔ�.*DF�k�1��֩��(Ղ؄ː�6M���Yu�E�2��5��=��N�6.���^R��73����	��kW�X�a=Bnկ?������\�s�ҕ,Á^��Lg
b#�C���`N�$3^��{J�].������I��(�aI�W<�nRLS��j�b�� �" ��R�f�{3�R߯PM��ݥ	U�������Vy�O�,pW����6=��ώ/H��Pvc�
+�'଎-\��s�T�@�Eǔ"��7SHF_�J�x�!/�H/Lgb�2q!�}jM�m���'�덼f8���a)�����|��	h��/�V��4�f���X��L;�Vއ���Z�ݔ
	,#�)�@ы]��<��;�8{{�q���B��^^�^["Y试�	,�H�&��_m�m҃@�,�� �����\�]�H���.�����vl����W8D|������R���d����mL�L��������z_�p� ��}�۹��CT��ח� e���i�� ��k�=]�����������\/H�\�p%���c���D�
F6{%DY� ՚������ I����͜���
m�Y�$3��f&����]��T�1դį�8�p���	��G)�Z�w�W���,�x>�&|��x�Л��\�߶���ϝZ��Jaͬ��v�G ���b�(XZ۔� �uр|�-Wi�P����m\��:�$S(�I���\�Q�����Cel�ÄY�F��{dº��>1�f�N++9�j��$�1�{xE&�R��U��s{\N|V \��=�>�:6u�3tW�'�[�P�T���(�d��V�'7�Xz�g��Y�|�D�DF�@.�����X���0�k��M�.�ff�����@�Nu
O$���3�#����!	~\Mo	V{a݆s�,����;b�&�L�1��1^��� ��)(��d��e�)���e~�/�8�$�R��nR��&l�� ��S�%�eH�k�9|�y��_*��BO����)��S��3۠��>�dk��I�Q���';�|���S���RR,��WY� #m@���9�yK��H'��v	�Y����*��e��޵G(�@f�ܑ۸�+��Aűp���oTǇ
����(f�Ib�
����"#����t����Q�P
�A7�x�;��r��#�b=\0�E�_����tT�x	e�K=Q1A���ff{��8�1x(���Zc������yh���ǋ�S4�(��A�+j? Z�ؑ�d�eG�7���ES���T�T�n<n.`^���a5����*a�b՟xw�Q�����:�N�ݽ�����E&�cw��7o?Y׸e-@v�s��r�&���{�"~�d�b�<Q����g�������*����5@V%����+ut�{/g�����9z5z�ŗ*C�O'�ۡ9Ϲw��+�Én~�?|I1��N��Sh�z�~c� NUǵQ�|R��ӟ������gNl*ڏ��E���oب�d\���d}���LM5���}v���p��D�p�٧���ㅑ����awe��)��xG��n�a��1~�G��Z}Su��Cq��g��ǩD��V��W�3{B�=��)_	�[�wa��M�� gm�׉����yX���j�����9�X#Y��������KF�E�t��x
��{(}Io���(tJ�c,�~�t�z!Y��qŠ�i��S4r�f���@�]��"���,Wn�+�/ϔÄ�7�Q�ɫMx���C��@n�U Ey���<LeN���E�R�B��MeG�����gwi����'��ރ�uw���W�"���*ʣ�6�[?"%����4I<v�y���K����
�Q�wq�
\�;�
��A7�hP��E���8���}�")�Zޠv�¨�b^��+M�g7��#�?�GT�K�yQI�u(:n��QT���t�����#�C��r�RxG��z�KA����KV�S5� Ư�;g5�����R��r��f�ɽ�'d�:R�TL��Io*Y�����Y��O��})C��dP�M�T���."`�ڬ&C28o;���uGW<�m��~�1�mh���{[T��z���Az��?*^�d4�X�bvL?����}X3����$��W&��+��S��x����0�L���N���f�J�#M�3g�Cr�X�̍�;M�CF�ǃ5�3�>G�=�����{�Û�R`/�0<܂l�3<����`չ���"�����f�'����|p�ѵ����y6�-K%&��?�>�~/.��k�h���N��X�a\*&ZMh����ݸL���V�8%u�Ь�E,B޲��E+4j^�݄�'���1�x̏_W��&U����`V^#�Z,4&U��<���r!Ӭ0h�6}v�2�PQ�42^hM"���(�nca��:��Z�\�}*�v�$�%{����l�aM���"\���Y���N�U=/y;Y5�6EI�E���6d;�2W��)y�m3{_%���`[�Jeė���9��Bs�5�2���ZrFz�����Z?B�FYN�2�g��xm���c����)s�ӪH�P4�e�"��e�
x��E�(",�!~@�>�SH�/�_�'Jw= �#F��+��-�H��V��u,�ǜ�X^_|�*_�̬-�?�m�� qx�/���^§�?��t8����+��,�i���$"�WJ����.�!q�@��;�T���W/?E�d?n��h���p�Ͽ�	N�7�;̪�,�~����Æ��[�����`����~5��\��ަq�ԁ�xz�F�|�|��x�����bb)HL 5-,�����p_�!�OH�yG�_�xh�;1�	0g����A5��X6���J���޾��1(��8�ƃ/~'�0"����H�ebL�[�QW��o���kk(`]FNԣ�J��f��hP�0L����(u]-��D>�EF���3�<���6�T���V���L����E��t?iAwc���նE �~�9���$x]s�[6�y^p�8��s"�G��Sd����q����	6���n�x,�o�R�G�	�N�X��.�0k�=�Q��!*\a*��<������C/�Ł p������MK{b���£�k�w��؝���*l)�)�%C63��E��PR���@��#��q�ֿ�$�����8z4��Og�:Z�y�J����YQfhH#C�7�^�IVA�T#����/-.�_��X�Ņ��O�ڞ�]E�ܝQp.�����骃�cڹ��윪cB�Խ٘n�x��Ԯ���?�h������N!V�>$�s��1_uM�@�J2Mu�y����p��'��̇�0�f��M�|�qG�%2��.���*����n�wt���_LY\��8�Ak�,?j��R�>g;�6v��;d'��K@\Pt�v9��׸��'��n�����C=�*��]ڎ�C�'�r���CDMx��jI�M��[㡐���	�c�?3�ޏ.�P!̘��8SLG_U7B� t���NRwO�a��)��5�q�z75V��E1YYT���ze�e�[���e�Q�[���]FY�6$�����V����E�f��Q�^�X���΄q11:�,ֱ�(+�u����5�֦����܌,�٥��8�=^�`ŏ��D��!�.�P˸���Q��o���Q�;���iD���Q��r�A�E�1�̠��벗��9��	��>���� @J��R������^�V ���+0t.���p}!���OEd�Ͱ������5N�G/	��jm�f�˲����;�F�M�6��C	{LS��L	)�L�=O�Ĺ5/�WȲ�K��v0H ژ��f�_����J��T֠%��I���k�S/�Y����-�8��oI��!��O��0��J��QN��=����i[_}�P�୘�}
-{�l�Xl��1��G�7�;�����(�^}�qQ+��.p��ʎ���["��r�R�gI~���Tۚ�g�d)���c�I��vi����>��h}��aS�.9�0��f�g�T�<#��ψ���d2N�����#I��6F1�2�g�,� ���LoG��h����&��n|����.xy^�#h����C�K"i�D�@yT�	 ���ӊ�ɹ�=�^�Q�����z���v�
���]�V����Zmf9Զ�e��I��2Ne��jh���=PY�~�<�Ae�j21�Ϸ����pR�Ԡ��a����ހSNl���M �[����M���H9��8���{;��[2C@�L�c���9N����ѹ[��\-/���tp?�eZP��)x�1�B,�V!@uЋ�j�U�b9w_��;�Ƴor�����U�G�,���{�]�z��wУT��/m+���N��_��U�@�&�ͪi%���W��t�A"r�-��N֞ �9銣��	��1��n�R�RA�q����V�ٿ?r�qPaa�$#7�ן$��ZH�u�+�(�v�x�E�w�1�� � ��2�f�\hQ���%��K�P=��
�y�@��7����7/�WR���%D��$]��C��N�\ͮ�i�k�6��	�wǘ��9A�`�Z:.��✎�t��Ǳ@	�a4Ը��Y���7U�d�^����OX�v��3�T'����$ �-�Z+�C�?��o]�)��s�dr�����&���n9�Q�??ĺ'�5L���E�K҄�mq�2�ezS�(�_hW`��8ܝű�Ek���2H��uT����و��S�>�$�it�v)o��.f��̕�o7���ѧ^�v��q݂5�a����_t��2ƛ�&(�D��eiDH.��ļ?'� �ʷ�M��J��x�aO
r��I63b�~��*�Ǫ�*	�N(0mlel���#p����	CD���i��\�+w%�b����E��D�^7�5��J8'�ꉺ�o5 ��~�*]��ےSe��xK
Mq<��Y��z��)<�/��Lѝѣ��m�Y}=�$ԫ ρ,_�6�KШ���_g���SE`��r/�Ũ�r�;f�TX�I�!�l��10��P�i�>!59S�j�E�ǹᑥ�C�5?C��)��·�h�'<�M�~?��	�P�l��c5��#C��寒Q�Ǆv�+�e�*�ֳ5D���v�T�+�q��Lo�}��	Zg���ӠvɒLf�=��kQ	F���8�s�uO�D�C��,%9���c��B߭�:+WKޛ(�`�/Oѡ��.�)=W��i)-ӈ��,v�?���g,P˞y���~��ޗА����"�^صJ-�Ӕ�|���ueg:F�8��#�5��D�����$r��=y;ݡ�Zl���X3@k�������������Psə�$6#�-�>t���
��$���on��ؿ��1-_j�+_�n?|��Q�U�eH�pS��N���y�6��r_��C��U%_aly���ڈX�q�Y�t��D+$D�1=��2\A\��}�� ��\A\��¡��&:�첉�#Dѥ�S*xVO��8,'�ò���x�20��+C��"xq#�v
�f�E�d�x�`�y"W�caV��9c�Ui�&�_��0�2��o�?1��'?]�2�7��ݦ9Mwe�k	�
iN�/ZʏJC~���a� ��pύr�Ȗ��;���5�
���n�\�	k�J�h��\-������	;?�8A	�FC}���n0BYׇ$Ŝ�������ص,6�C�]�s�Xp��9���l\��"@i�a:)���@1'���=����M����ӿ���D�n�t��,�s��p�q�Xllȭ��;-d�i@8���f^��<��̾����7�BǂiT� %6:��s7� s^RfB�4i拝��26ˈ��{���5U��i����)F���Ŧo: ���+Ԇ��:���ن8�Аk�	�	��u���)g2�A�f��K���{6���34��Z��5�&�[:��s��	��2�,������[	B'�6[|����V(_���3]�خK�~N��f��՚m�U�j�:����|���� �)�P�Pɉ�[�F��H�8c��8�ٜƥ�kU�V�d����EC�(�ƹ{¤�M��A�T����Oք���S͵� o�%�R��C{|�V����j+�Oӳ���m�f3 �Tl�m����s�P4i�����	_t`��.��dBÞ-;��
�Fɓ9U秱{��1�]�����k� JQ��0�����8�P�Q�D^��T�Q$Nap�mҒE��!˄Nh7��>GC@H`���l[x��|��V�W�� KZ���0q��|#���δ���yL'��6�-��7V0�����1������@��~�݊�8%����WM��T�*y�u��&$/-�DOi8�/d9�&¬.���E��E��CIÊ,͐���y��
�.�-���^3,�@��?!)�Q$����I<����ٴ�sPH_9.>Z>Hw�'�`Y6
 ً�q�Mp�V-�.^ʂ:o0�z�%�C��[���p�]x���uYzx��k����mU��K��� ���
f��~���8a��@;�^��ϧ��P���u�l l�����ߠ�W9�V�!u���,��n��j��2<���dvJY}���w�e�TyM(2#`�ec՝�	��[���!�������p..�9��.�OlUc��q]m�����y�1�����*�H3���[��H�7F�|�K:E2�`���hC_�ӆk�.A͵�I7�xrVu�zh��{�d����� ����O�r��y�^������d�SM�?<�c��������,�A��"ݡȶM΍s)x�
44�R+B���x�nM�%�Ew��[Wn=��ۀ�R�<���0�xNJM�Ĉ����	�/q�b��~T�ϊt�Q��hN����W��6z�i��5�S�����L.�ſ �Q{�{_�{�&	�Ƿ����8ף���$iH8n)Q����f��.G�G�h[�1щ4�{�z�"*�K�	�'Y��Ov���*�T�:b`M"� p����Q�V� Y�)���>K4���kG�Fq�A��������$SH"(��c���˱��	���t�f{E��N�h�u��c��8FG������e>�rʂf[v����>�:�	)�}*�Xd~��싑R���ͤM��1����V)�ʐ��ta�(����B�K����RP��%�',�`��PŠGzҮ����cx.
�;��*/����~,JWX�e+�S�G�A��B�x��;N)�,O�!�����1o��~�G�[w�Bn�Z����D����-��8�U9Kl�d㮾i��l�c��B4�}��K���ꔇ�-���m��������J�@�F$mȶ�}�p�P�޵n#D��hЙy[ڕ���ǻW/]��c�^ٶ��..wZgygq��¨�z��,��M�BM�����s��ѯ��Rg�t���/�������pH:�������,����9=K�2�2U��VD��a�L��udg
�f ̼�W��܋�#��L�/��ư9�Ji�'e�����W#�drø��Rd�v٦�*��!��M��k=�I�a�v���7é�~}>fH"�!�?>/��䭨��ZN��n�%�,)/�(�����e㦌���A���	胀UbRŕ��V��`��:� 0]ɮ�I9�YC�_]%nc7��s�� �(���l���t���Ȗ�D'RI�ս^�F�$�.n'���K/u�7 �z�nwK�ß�ʖҲ�0%`\��䩇 6յ����x�ߞ_
���l���pw2\}�Y&��C�l/W�����|�="��ɤ:�2l�p���ˤY��������I�j���hkU3�Iw��_�I��T���z�S}�/������I�����m��K/��Y%���l�ʗ5����<�o��n:�rA��0p�r����$͛�=�H��R��-���J���6����~3�����j�d���I}��v��)a��1��ͱLF,��>p	�PFf���:��%\�-|)���Y��Đ��]�j��a�k����Ud:~̔+�=e��I��0z)7����5��\��9<L_�M��
�&��uG7e�͗b%������C�V������a<��(l.9���hk�k�T��8�Ƃ�7�IM��l2MחM��58t��'�q_s�.�����:�*+]���;ujW�9�1L��M�.T�]�d�w	7��P�vZ<��#M�{6��x̓��w�Ee��@�{�@��E��C?��˨�Qv���OX���K{E��2O-&�-/Rš�;ѧ��W���}�jW�ꭁ��p�� -9��͊�2k�������٬�_�X�O�Ei{� j�S��r�{ �_5�4���Z�˞jlSˍ aX/��.R��
�]���=�_I��������Ag�*MB���Y�J�!����>�X��@���!)�a���9���sD:Q�-VD[���b������r�g.����	�x,����qfU���FS�������t#m�5)טe�f��eY.��Q�q�y+M%o��A�:�5v���
}{G���To.ޥCF�Ğ�D	_�@��>�D�]|i� �N��,��{�kԞ��J>A껃�LPgu\���.@;�]���!V�WG$\�E�����P�Ӓ��{l��/�=�O����#I���D9�b�\c:�B�Z=����yJ�2���k�#F�~�'	-K��jD�F)���{/\V5i&Z|�v�7\RE[ݞ��)��0�8X4�'k�<yssu'�xNQ������0ϵ�b��2(4xy��]&Y�&��q�^
�++�S������̱�4��?j�,�<3_����s��Y� u|�5_�ғq\��s�^�y�"N�T����מ+.Lm�j�8r^�<��
�<�<��'�-,,T��4���* �c�������`��F_���*B�.����LdN�s���e�$�0�5?g__�A����!/y��L1�d."�z����$�`�����bR:v�=��bLy���o����%T���lb'��Z~���>�,%�t}65�+oCÚ��j��C2�O�X �o=��<��MfI�.��Pt���Ї��F]`|�V]������@7�lc�����4���A�x��տOcAHha2%9f庞�9Ҭ�����6U ��%���D&sw�SwM9t
�]�X,2�1lp��f����k]�)��-��!��b,��&�F �M�ba)W�bs�1h+����:��*���ה�����rs6d�?x��pKۿ�T;���r����Xa;���2�IN������p�Q��4c��[q����s�������7��z��k����8��񾗣�`�;z���7UcVɶ
S񾿕ۡ��y����T�ɥ��]�Z=i�N1�U.�h[fmj����w�X�Z|хIB[�`����R`)��F�g��)2���(���"I^�cPK�퓁�~�4P�{����C$5 !� a�o�|��t0$�Cq?� �v�lV�%�=h*9��������34��uXأ@�d�D����֞�����cxV���g���l�����G�r�Q-CGƪ5a��X2.QN{��)�sA�%��@5���Q��śQ
L�A�� �<H�?�E$��qyT~��y�0Z��T�6�1���Z�lh��`�h�²B���F:�U?�o����q��\��F�&JG�G�Ve�f��n��_ѹ�句R���v�pX�Vq��*?��9�L�i(o3(l�9z@P�D����j-�q�Ҋ5	�h�Y���+���SoDc��|���њ�9����:�A��Z I	 �����8]{ ��J�gG�J�f�ʷ�;��� ٣���]�Tɾw�n⤽�s�I@�BT|�20�'��Y95��/�+[���sJ�]bUa�*��J�ۘ>�V^����V�+�E["�����h~?9����a~1�JvM;nl��P��nW(���dR�֠�@�|'�i�`��L� ��%1v��S����O��6��^:��Е�G�4�0$�Z�-_4����^�ⅆ�¨��6y Ų���U^��O!�З-�X�Į�J=��'e,���Mz����1S�9#X���MM!���M�Ӿ~�'(jf��A��@2����Il�V�TI����΂�^���8�/WAB�]/ �r��R��+�WDR*�)��|H�ݮ�K�%���	��ao��}с����jW�v�Ů���5_�;��-�+�wg�>/$P𩳝�J�켍���}_%N�?���+��@{�s�s
���J���m��se�D(�o��׬	��bf�@_-
�����3����,�\'@���0��|������{9M,��c�?*Ɣ/=i5=u��>	Zߵ�h7������Wn�	��T�����r��3��'�Jp��g.L{I��!�~��m��)m�\0�T�`��<͌��VG%�Z���Cq��--���E#�{���<�q�
��p����`��Y�L�D-�Q��fz	O�ӝD!{����k��M�N*��I}lP.���oR�r��a�CJ�b�6S���:{��`PVy�1��S?ىm��V�):&��L\�]B=ZV���ZsG�c�%Y�&n�U��؊:t���N=�7��R��&���A�x��D�@�|��nۢ3�n�S�3ܪcR)�ȭ�Օ�?hL�{�}a����aj�H�^�k����ǯ�F��e����ϰ���1��W6I���[�[�k�oM�{q�#,-�{�Ơ���3�_��C2>���&�-�� �3���8�&���cau�|�R��1�瓭���lF%@����E~�l��������1{�v7��d�ZWJ�3��_����MaoFtH�R:�W׉ph��m�A����1N���-z�bM��~�>;
�Ι�#�6U"ʴ���X4Npsa��5���,���(*�$Zu���iS�;t�>4A����QQ���{�d�(p���D�
`Kk�蒫�v`NHg,f�wA�PQ��(�[H�$�x���[ځʫ��2�{z_�*y	D :�i�<�W� �ڮ��lT9�CU��3Q`��
9)F7���q�2Bw9�=�|�5p�D|f��l2�μ@��i �P��C�̶�"��sH���g��nm6�e�/ử�m�8Ñ*[�MO��t��_��Hs�C�?�(a.BQ��ꪻi�B�<4̜g*��zd|����qP*�pg'��Jcz;�N��r^�i&Y��̢�fE��rn��UfZl͛�;�=���r�u�R�#�is�>N>w�d���y5(RkWkD����l���\�Bn�W���ϾT�4�=�Ya�߈%���m�:�����fu&d�w	M��+�SwЫL����׺
�������Yv/t��(%�/ ��/ն���e���(���c�c� ���op&��Q,�H�1_@����DK[�J	jP����<��f_��6��n�Blu������d?��@���(|ɖ�j܀��-�w����������rB�YFC�Ԛg�.3Z�����w^1EN �N���P#6R4�Q��q�I��lI�v���u�����SZ�b}�ܚ�B��[i�Z�zZx˭��r��~X��5��h�c�m�n�oh�,�
�7q;2�hҡ��2���XW��S�Wt�E��M�1.&�M2�AB;F� *U�jx?�j�5iåbņ3k�W���9}��F�Y�b�
 �z�>v̄JFLx
%ODF8�g j��	$����Oal��|�i�#z���t��ȡ_�}eݟ�!��� h"E��DFN^�kM*��!(�"��o_b�#�����Qڇ`�E�]bM��%E���1���z��i�����A(3�8��������?؈�e_|J���FSR;�X��d��H�GY�P����!�ʣ�:�e��Z��po�������6���'�bE(-<�e�Hv�O&�}�W��XLn������#'9ħ�k�'�5����M���ЇM�m�!�;� ��}(y��3���Ȉ�� t�@1]$9���B�,M�]�e�w":\�]<m��fh�Zx��JB�2<� ���m�)5T2=���v_&�"rf*�\zÛ|ڰ�So�
�B
&�s�d��u�d<ň��-k~�4}��}�L(P���A�hޙ���<Y�U�^@�o�@�z�a̞�o9K��cFk(:q���҅*�n��^�2��^.�ՙe/�r��F�t+���3b��E�����������:������D���6v'j�,V�[�a*�:pb�3/wL<X���w(\�/�"�07͎�	:�y'�!���ύd��(�&B@�Lm��6,���J�p{_�}b�'`�D`�mɐ���Z�ワ/�߀b��AQ��b��n���hL�,��eow���b�i8�g���C"���]G�0Dc�6_TKL�糘,�>���/�}sT%
��'"/��պ�g?.t�������;U`�aPx��̧]!9iƞ̫v�	���x�|8�R�N48K-0�	<R0�\�渶�1�x�B��޲L��(��0����Bg�:�H�^P�GB��-�f��]�S�cl��3�w���`���` ����aT��� �_!��GZ�eD�u��V"�NCA3�>3��%������jw��U�y\��͕~8����F��<�
����,D2��^�ǁUH�:�%�f�Ud�"�V��)жd����[{��ʅ�����El��] ;U���VZ��Ӹ)����K���������Ny0�hM�2�iT:+O��{�
���m@�
#�jv������=��H��sO��EN�B��OѺQ�/�E?�c2�Ęf�����Z@�xF2�Y�-�Ntf@3ӫ�2��q@x�ӝ +�.�e�1m\��?^*#z�@OD�c8�"��N��z!v��&��%����.��M��ÊP�ɀ屰��	_�(�Ÿ�yd¶>L�#�ԫc.1�����0�)f��KWF.c���&��J:8�`$�4�5,8�/�]�7T� ��&,i+-Q��F������N&�W���Z��R8�oDQ��+�S�'�[D��à^��}��BW����E&{�ifL�-Rv��K�y�C��⬌">�܍J�?>�h���h�:3�h'�ꏭ��_��U�
$�< ��@G��sj��uBJ�q&��x��}T�ZS��b�p^���$'�����Y��m�o'�&gˀmm�r�����	��G����kܵo�ȵ�.�ڪ"�٤��l��I�u��Te�B2���r� ��g�4��"�L��9:����hG��FfM�ߕ��6d;��r��ǆOt~]<VG�R������R�#8h{p7.S����q��I� ����,,Y����"+<,���⟚�����PP�u
um'��.��_X�4 ͱK���^&5cՁla�]����1u�Ţ��SO��q������r�������c� �<���D�}�'z��×�L![�t��mT���ɵ��rǼ@���� ��\M���LѸ�x�[��v��?�Ľ)������y��4G������Z|u&���������:�'d��p��BPqqD���|��� ��*���&���+2J2��*���s���i��x�[��B��cz��ji­%�Q��������L^=>_��x��%�V0ð��N	4�+�E���p!��(�![ɻ���p�T���^�Y7�*{=��P�w��� �3��[�qr�P.�蜰��&���N���0a 6��M'���Zf�����Ah������JF�l��ԩ̖h��%����:)�/=�테w�m֛��r}�V
OJ�� .q
��Q�_��˚rz4`�����M�T@]<Z��k~Z����O{�?�Z.R�?c�����4�Y��G�j�LH��0���c�ˀ������S�2g�9��eԴ�0D�"�0��]���b���4�4["A��Ze&��2J� �4�ɀ�"���h(}�:�f�î�iր�M���@�2���_Y�W��{�i̊O��n��w�nY�#��2]�����ُ���ʔ��.P�F��048��-D���5%��7�`1�|x1rd�L!�['�F��-�#������ۑy�7P>^BWH�@�i�b�Z���x�eC
�F%���.�WԴ�Q�[ {'
��	�N�Q����fE+�����>n>�F�م��BTl���ə�},��o���Ϸ�V�*�E���s��"FmY,�A�9d8;�T��!�*g{�Nn�I[����t�Ő�"%@�E�Sr�f�2�=��4�����D�=�5U4��[��P�˿����)M�?&0���ۆ�T�y9���J�N��Ҍ�濠��h�T�ױ�>'C��N�^n�F$L	$r��� C/���)3{ۦ�i�
�xn`�ı||#k'1Syε4Dp��*r54��s��"t��eu�D�K�ȈB**Z���&�H�L�3���Gh�BE�M>�u�y�sן���Ԡ�j��rɁ j�B<��_��B�V}a��Lي%��qM��W^��\� �pF4��	�������yͭ^p�q\?�!	; =R�o��|G��7����:��$0��� |�ƞ�����ߑ0�V��N�"b��A���\[C��1���+��!�;�a.�I��5oP����`�G��x��Q3ń�6N���6��4}U�-K �oR�R
@x]H��1oD"o��Hi��l~r�p�9,'ҿ�9�E��E���.�MY���q���ܲ-�h����I�0���mG��{`��Z^�R*�!��ON;�-�狥n�s�����0bby;>��;nP-���ô=]��3n
A[��U�L��0�N�룟��V�������e���_�d_��Y ͼ\D�b���1��H�j�õ(4���Z�ܺ��&B�t�[��(��w(�	����:$S�0�3ٲh����9��ǐk��)y뚙�t����դ#� ]p����u����y�Ԓv;�n��y� R��.�i�H�=�ٍD�o�=b1sp�02O�D��86�6���6|�+��%��C⪎�'Z�ڛZL�X����<!�(��gE��T�'���L�9<�W��U�cR��t�@'BȊ\��7G�YO��_��S����@z(Y*��>��%b':H�訍j�1?�v3�83��bq7v�#?���:%`��J���',�p�vO���EI������ґ��O\�b'�m��1�'i��:p�y�B�	~e�P���q�T��t�Ӫc� �p�������~W��!�O� �^hZRI�|]xYLx����8j�����zo �F}��xoT_(CyF����H�Lj�Ny���3bb=�?z��`K��hnǩq=���?[H���e2Xq�J�r4�K��Sݑ��d� ���1����&�;U�v�ns��*�����m�uT%�������� �NU�H�g�M[�~g�m�<��!����o'Ʃ0��4.�ˍ�����DA�2�#�`��r����H̯��:����0�E?�-?�|��'y�����J|˨��9�6��~c�H�y!D�D�YRy=��/kXTJ�|����È:i��[$a���M�|�{�_L=�'(�F��Nv2cg�����icQ�>�BίAx��l~h.,���ɚ��IZL+�z�������AܟPZ's)��^���C�V���M��>�Ri�����@��q[$�^o���3�-mY1N���m~3��2yw�ҩq��,M��&f�@P��H�Q(���xWB��aS�&ONx2qU?1��@j��*�Q�_�"�&S�޻��CX	��]��!D�Zq�#�2����P��
 |�)m�+k�%���ٜ���s����i$��x��)�`�jY����.YᧆY�2c�GӅ������ӀI�	>�0�r���M��7yg�\����w���Ӣ�u M��0�kP�H\1�
��"��ap=4�P<��@��N4u��j�'�x���Q�C��m�|dY0���ŕ�@ $1+�l���k��Ѡ��%���
�����V� ��F�F|h�#�޵�c��WZG'I�|T���El�<w�+�w�/��ʝ����Q5�h�"�8��٥���t�Ӏ���d��f�$������Ml��	�`lb�@��J^�%�~E��V�^�*L<�'k-0��/\��Π�&R�kR�bpoO�1Ҝ��Y#A�%�^.v��PG]�WZ�NR�I�t�9tU)�~n��~mL�f0�wWE��禱j�}mS���xEX�˯/����������o%�����#'X�F��!핓Z��&u��(Oe:(��叙�oW/�����s*��y�b+���7П��Ns엲5Cfme �*N2|�u#1�"��uH�=�Ʃ��:��^],v�~��5p&�)"��zS�B�oD�{�YÎͺ����J��H�.& LM�yt���	�P��ߠٲ�� ŧ�I1��:�W�oJ�Fcf�2X��AN=���C7_�� �<㫄����`<ųX9���7Q�'�ӢB��DfØ�~+��������� U��aK?�ִE��y1Qx���z�
��O�>N#M �¡!�{
T���-���%8퇂�X���'n�����\^o��I��sG�%�{A"!�puB��ʈ�������Z���Ĕ��a�L��K�0��K��f)�!T��oE�?PT� 6�v�C�;̆5�XӈTb�'�io��C(�9ɳyH�u�+�fc����V/�`�Ǥ���y>vδ��g�ՒP�%�$QP�x3-���[������&��)��S)���R��g�qt~c�Sl���Io�.IbW�ruw_\�J'�Gr�g9+#o����=��X�����5i2i��ɓ-3ʽ)���I���Q	����r�N�h� ܙX~��ws����̛a0�MP�x��;4Q���"�~�r�Rw������$fh�ڳ/�i����@Q?�v�]zf0Rv�as��-�O�_�d�5�>+Nc�ė+!��Ԣ�m��,�ӻ������������햳���r��# ��)�D�w>�V�A�nh������atx2���/H��V���5����P�*-D��� �X�k�G��d���t�iP`,���`Hcj��������������r�]`�@6\����>ERO�i�wtWL�/�/X���]�1�"���x_e� ����2�4gb�p�+��q���ɞ��-ɶF]��ϡ��F��dsVB��GH;i����`c���lc���\TsX�^���zF8�.~!����7��D�vpJ�<�@����?G6�uX:���|ib��њ��9�����y|1�]�ә$���t3*�O�������@��C}I�G?���Z�(��]��.��!����[%-�������|U&h��e��H���v�(w�7lk�<���"$��!�?�H3�y~e���,�
��}0�� ��� 2���a�����y�~����)$"������qH�f���e��0�'���|���e�@,@��1l���x��N��JW���)A�����@���ܒ�մC}���U5=�r�T�@�*{�r��6�����XV�@�X�Bq�o�sgF�J#���A)�l�����;p&qn��j��jR�ӰV�s�z"u6Ã3���{�8gI�F�
d�oxy�@rcGT���_|��V��ߎrN���@�nl^����(���C3��y�0��g@���e"�*��e[Z�8�Bɾ�I�����_`��j	��@9B�һl��G�$��5.�-�qb���P�����@@-�	��G��W|�H�?ʃ<�tg"�N�sw���84�.*�UF��^%������aך��n�n�\�i�H��$�	�r&��¿<�<+��@�%���Fm�i�B\�A�-sa�f�/]����\�	]�ɐ�N�
3��b�XW��{��X��&�(	�)�3SP�(�p�g?��b.�K��6�FY'���Ui a
������ڮ�JW�4@���%��(g�j.�l�c���������I�E���x�[uE���A��)�cr��Ca���Ȉ+�=֐��[�A��emXJG�CQ+�����������-J/a��v�I��4p��X���F��e�4�ujm�U�}��G���&�dZ��[�˻~r�|��O��+�X|�a�3[~3-{@���#���23�L�u��/�˳��K��{j�/��˜8�BdZ�C���	"�)�oBڰ�{��h��W�Ź�^�?�#�j��;S��{o� �Z�D�'�LFV�l�-s�C�}�q���0���W�ǰ����UR���ڳ���1Sj��4�	�V��K{�z�:���U�_��qd��^���t!��sa�:^�{0�Ң�Ot�Q"��mU����4�I^�xg�v���ĩiG
~v�o�1v����rí�_�+k��?+��O�
\��Q���a�xG� ���e9�߲���~l��u���䍔<�^�q�(=]j���_����ޕ�=����JO�B�Ҭe���#ﶙ`X�pV�@L�UcҦ���ث
vOb��S#y��=�!���9����\�������"
E�R��(��ě�bz
*��l>�:��Oگ�{eN�"SF+ɈM�y�,ٷ5R��?ڏ��g�ի%'T��xJ�Gt��	��6�Z��q�a�>������y;��k|	*#pr���Jd-g�%.����;/N�m���.X�@:�$�*\[����x����:��;�n��X��R:�P2�f�XYI���s���z����s��~�X��I�^�&�~�K�⧴��+<R ��+��9��
�u�LA&uSOǣ���1ܷ)��{�YRF� )x-�3驱��[��|f��҆�%7�_�ΑD󎜒@}��k�~�C�%i����C��������~Ҁ�,�Ot����0~���Py�S�e���g��,{D�F��/JMT/���Ѩ�uug<b�K�f6
ԧ
qkN����\?n;m���}�m~.^7��Sw������9r쐧�}V�t������a!�4wz& oȏ���T��)��֢�O
�{��J%�+��p�����"\��4�����,�mWS-=�H�2c}���x�Z�3�g+bgn�Lb�Ɔ*�Ƽ�0�v`����J~��������^;i����}�T��9�D\��,�m�n#�"��G�6L�b`ˢn�J��a�
*j$ډo��S�AZ�	�&Cq��Z���ڸ/�m@h�O�'^�z�"e�QH@����Hk7Q��w����	�:�A��=m��(�a�DTIw��.�;)���i��V��e�GtM���S#�iT�m 7���$67�˃� LG��;N�?t���a�[v�������JSQ6�������H�+Q�p[����z>q��=��%�G��4+k�Ә���g���\���/]cƁ��u'\"}��/Ac�t�ݴn�ǩ��>S*K9�eL�8�qM��7�A����8ʽ'͛j�QL�/|Xw�.���!-0,�?�#�EUZ�+O�=hc��c);�cb$��^��o�����;>`Rj#b�Yo F〉��'�y�T��K
F��F)a�*���6���t���$�H҂�,4�U�L�݊ˠ7�l��q�OXzF���ǡ$ ��A�b�w d�R�oW>$|���0��>����6A�́L#F������К��f�&�:I��+���e1#@o����e�=2ՑXM�)�7Uy��c��D�/�*�ȶ�-�� �
X=�c�� d <�n�d�)z$ܩU~0�-�/9�f?�a
�s��9dzsؼ{�EA ��4O�X��Q�=�{��6[k�&�A�G��n;���=��׽�d9�,���?�� /��\�HZ���_�J#�X�u0�������#y�*���*�\�$	&b�-A�Irs�<[>���9J"�&]/TH�����Q�f5hx���U�>��P��Vd�9t$�^򨌉�4*oU^L���z �Կ�+g�T��m̒t�?�87X�H��?�DU�G��X̏�j�����|W����$tcs�%{�_[���ML �r�6�E�hm�=Oa9��Y�]@0~�ޡ�/،+�=r��8�"�IBh�ay�`���54�gC�0��H�'̓����z���2���C���	�Z��>�)�4ZM�����ր�7�k<����E�paL!X�(�А����2rq%��b�Y����;��9SO�G�©	��f���Sa��ߡާ3�!Ï̱m&)��KVl���~���ڵ��F)�5���c�c�����#Ǐ027���fW�&tD[n,ۼ�������w�!�޺�F����=ԙÉ$�t��v�j������?����	 ��9�R5;���LR]�ku�Q�my��8	?�/�W>!8廫ǜh�R8�V�a��� �63�=�A>g96T;￢G�m{�/Zي�eJ'��_ǘ��
��HNj"^Oߘ���%�5�\����m�'�����b[�bEn��8B^��5��B�&R��,?6�^�L��I���Q���?�N�@��D���2��H��H?c�>��~�<�����W(Z�?>/�^_;��E\m5n�hX � ֆ���>Q��}�V�-Q�}��� ������-hWǵ�]����"_�n�c4k�k�Z�vO�H`�TC�_4��V /&��@}s��s�D+��M	ĳu�~NU�,�����x)�͢��2�!���Z�+/!k0��W�

��Tk��C�z��/�G���jm`�;5�#�Ǳ���Y�7-<�Vdˈ���;��j@���	:��f;C$U*�4r�C��� p�o
����smo��v���&�b��k(�e�M;���~Pc�n'�U�w������v�,yH M��n�u��z� аjH���,���d)�A��Sޜz~�Ϝ�,��K�ؗ�O�#�L�;V��6������~qrq�>'k����]����˽J��?�}�eT�H�$���!GEar��l;?o+��nL�|�8����37�o7B�����MDX��j3W��V�1�O]�6?>8�3W��Ds���{9����nD�3���E�],ra��?������ׅ3&�ˮ{r`PX���C�Ʌܩ9J0*��o�q���J��p�K��ȕf|����-�WO�rf�Q]~+?*�J��NW�!����T���%�C�d�´��~��	!'>p&!LF='���D�u?��X�B���n��"���:�8�g��H@,/�1N�(R�����I���Kb�΍�=�+�<����x�ۇ�?�9�Kʞ���[��M��+�>��S'pً&��~�0E�*+�V��<.��X��XNQ����K�=w�`˾A�9f�9�J���n��2�-\��G���&�217�*m�1�!�m�8��<�PT�'��ǐ�����<�4[/"�r���(���M1MG�˄���Ǣ�}ld=��$�,��W3�t�O�3A�	�O�nz���N���ׄ�x�pjč�_(.�^#�����؎��Z
Zp��Ұ��N������l"Z\������X�A���	�4�W�"��KC�)I�su ;�I�ρ��l�{(ܐ:6_B|�Faɻ4}_��;��R��*O�`��V�o��roˠ�Β����F�e���INs�?¦�n�N�	I�w)�AT�fW�w�D����c�"<0���	7�Y��Ԯ$���LE6���0�<b9.S���C��&g�_.ĭ�v%g<}ǵEh��k��'Z� er�:�IF��F�d�U6$� �f	~�ֆ`N��0�a�����&ٛ4� � �����JO�Ɠ���e�'wO�[�R&rj���5k�
^���n4�8J�_�|A>��nc����%��zD;̶��n��W< ^*�P����k��M��O-������'Փ;�Z�1[�l�o ι�5ǧv���N��KqM'�!�������n��/���7���+v1/��w�� �i��%z �ȴ�},��퐘����GZ?	�`(���sdZ�8*˫a��A�E�v��+<�c�'5�P��M��WG_�}'���Gd�T�,BE���1��
�b����W�������[��Pf��9��<��d�q��vr�k�a+ؤ�"S��]h%���j��ƶ
x4y7�������n�Cj[�B�C;�����}�{Y,��Ps�q8�����ׄ|��mBOB�dʷU>��� ��P���½�/�B�!j*B�}aW}WV$_��0��H�2�����y��C�t���e���Y�(�|�;�Z��
���(��B9T*^��|}v^�8���缢�������p�3%`�,��y��ˑ[�E���_*�%��d��rã�U�Ӷm�[y�P�L���r���7[����_(_wZ�m�W%.u�x�Y�_�ZNJ��->�����B����x53�1�G.��X.�opw庍Io��]��#n�c6��8�2�Jjc�np�0�<��VM��C�nL�_Uz����i�����?'>d�u����L��<s�5��h��z�
5!K3ݽתm��-�
F�l�z}�1�� Q�?��襙.bMD�KS �[�Q%胍)��KEn)6v����E�6�����(�8���������Wg�7�/�X�u'��b� G|��=�Z���>O*N"�^@י>�	�z
���Hb�B�H�*��ܽL��}�\]�(^���B��5�͊��É2>�9�f}ܮ������k൸�i՟}�mo�k�]s|�Zzl��蠺�_o^WL[نͭ)V���<���c�3T;{f�r��D���]�A{��M��f��N���Y��ٌ�B�Z`�3�V6��!��ă0�a�L�� �A⍳��I���o�"֙�ߛP������WE���[LK
V[8
�<I,��U~����"���b��Կ��=�"V���b<-}�~sb|�T��EeõKq�ޙqB�Y{;ޱ�a����H.�q�.�Ü�VB�p���Y��+ix-|�W�cS"���z{@��o���G�������V�#��~N��9_����E+�\0��Q�CIP��n�_�,+��;u,��/ԉ�j2�O�9���:��I7�K^%7k��^)� �cd+=��/�������恬U��-���G���r�(x �rK�1|f	9�Dx�y�=�6�!�V�7��� S�+kX�۶8r��XW��D��3�j�[m���eA���_����_D#	w[6r������m����V;���ϓ��J���c�V�	,�ӄ g{���MRY\�SE!~B���4��ܻ�Nu��.���G���j��0��A���;�!�NȔi���R��{I׮�Ǿ��=;��!�vD�Dq��h�b���Vm<�7���ςv7��B:GR����$���ebV�z_����.Cq��h�upS~���4q���Ts�`dO�6'���i.�
q\�j�!�.(�� ��`-S?����/�U�9pُS�E��
��jF@��1�6��i�6�[�ᷕ��O�-˃�;������%�>����H&�:���Sñ���g�n����#��0 F'�>���61q-�-e0��1��M߃Q�y2��i����9V�b@��^9����@3��دS1}f���*�'^޵N���QseFN{�#s8e����{���MJJ�XjRv$�(���*ыC�	���x���C=�w2�g��& Ϙ�sjzY��B۴��#Z�o�υ5s'3M���:;��M���� e��Xl?��z��	���v��^�*P�S�c*�-�n�3��5�k��Eߡ\���n�� +<FS�f����v�7;���5Pk\/���IG0���:o�G~�x�+�O����Ȫzۄ}n��+��BI�9��s�ţ��}�Q���W�[�^�2=����y�_�i$�}�lJjIZ��M0S; ��!Лz�0��h䟛�n�_�Rb��~�,�W\�M�������Ct89�����ByP�x�z�Ð�3�?�I�Cz8#�`?=�9��n累:`L��ħ�9{�̐�'�E�"��덧hA���B�#��Ed6�Ŷ_j�֩L�A5�k����D�,qԭ^�,��%��$���ǧ����滤�D�y�A��>ƝN�;V�.!nm��M�R�Y
�ڥ�������-�(�2��\dr�(x�h�h�m�>���iv������ՙ�D�v��	_F�v�t唿4�xs���v󎏍%�O ޤE�<��LI2R8��}�l���n�iU���q����|_���^=���pС5�z�1!������z�ȦW��}�"��/�ʟ�j�8"-��� |U���KB
�y%�:�O���t+#4��L!�����BCZ[������w�R�.~�J�C"1�ӑ8��^��zD��R�,�q.^ 6[6ĩ<+sިٷ�1�2��n��8��FQaȏ�h�!�Ѥ#L�izo8�e��mӰ�b-ԅ�q �;�y�yyn��M�[��`Q��L��8Ua��/J���8�#��^-m7_}n�����a�Kv0�{@3w�Yהq�M�5,��#_FY�-�J^D	xv����E���o�����兞M�K����A�պ#KG!���w���.��Zx]�]��H+���t�}>#W�v�����P�7����A��E�j/C�J�
�g[x*����i�Yݺ·��#���
�A�,_)\�:�� $�Y�uՆ�s�s�r��zi�P�f Ғ�Hh��-�+��R�rٟD�H�N������e/�2�禽@Tێ)���&cE� tǤX�P>Z��Ȁ��1��!� ���r��@���n}Έ!$s���*�ۊ��̫˦p�١�:|Ѹ���Ygz���<�]��v9��p�'�������BZ�X�u��:(&�b���5Ŀ=]��Fyï+2'���T�^�k��PL�2�VX��yYc/ [1a��gq0�i�|5jO�s���O�-��\���!�.�
x-�n>����Ih��V]����܃���;M��2n|��񙻬a�$GG�G��پ|{߻�vXMn�p��d�!b��;Qi>�r;�;۟1ce�@��.>/tZ��I�7�K[�K��F	G�ia�k$��V*7���"]�W���g֨}��f���(]���e���h)��%��r��a���=�1K�X=��V-Z�N�+����I���&�a#01�*I.�gX=��"�dA�߼Do�CI7&u�܇�@y �]#�fU�ԍH0�׬~������e7Z���W7��E�X2�sTI$q��edh�(��˘�����v#��
��9a��3y]�����fWTk-�F���\z�7��"2Fɬ�A��x��&��Km��B2��� H?�7�;O�K�J뵶b�w��U?��4���E(����:�jM��\^��Ca�Ǝ���0��f�y3��M܎D�>�S���@[�|�BM ��*j�yfge"���jX��Y��LQ���f.pb�2~����`J2%�����uv�e�w��ǹ����;�Ɂ@�}X���@��.���M��F�Y�t}n����MoZ�Ҕ�`�C�ҁ�Y�暪e��=d2����e�T1,/@�(c=d--�c?�6emA�^�y��
+���!�6���v�қ��S��F��Od�}���SL�d�S�i+�5g2џ��c�{cb�������t��5��*�c:׿:B���h�b�Á�0l�z�^,��ZKE��uyn2?=	Kq,�Km�%g�����-��RGm@a3�p����? ��l��"��L��K*Dje3�p���<�/A��5,��S��7$�V"ZI@�_I�[IO$�O'#]�X���e�W �r��{p�ɞ�z$���''�HPE6�K-;����<������񗟑��V,�H���x�	��]8J!m����5�9�ҟ�T=p\���w�'nT���{��!����vjusg���J/|�������p�<ʷ]�6��)66�<��`����O���0��s�6.���$��pګ�y�'�!]&[�<��"�H����c]����ñr5�e2���*�a}pYUٙ<[����6(G�Hɰ�v����<���ȸ����h�c����wz��;u�c|���҄4��,�e���=.���X@^dww�?'�1 g�6	@H�`k7m�ݖ-��g҆7�c��T*q~�.T�*��^��@BO��L��E`Ҏ�\����sc/���'$�ε5~���oa�etF�ڍ	��v>9�>7��y:�$��(iL���
䡽����Teƭ��8�%��0!�h����&嚍�κ�p񬹘Ǆ�5�b|ͪ��\_��W� Ms���d��$C�@+�½	��$Ǽ���D�S�]Q�ьr�g1�L-��j#��I�ƺ��[k�GC\X��R�˅:ԋ�H��,�w<v�ˉ�F�-� hp��n��T5��gOH2�5�z�k%B���~'�F�D��q7��{�Ƅ�͹��y�b�Cd1#|I�!j��F�#o@ؕ½�Mm$������nT���t�B�}��p�ך*�nV��	�q��%����k�&�*kN���n`�A���� S۽��%�!<�{���Z����CZS�01���#�}��&b��p~��k��4u��6��F��KQ<�w�� t�:�m��U]���6��ri�`T���d_�Ě]��P�ֶ�,�7[�6���=8֬17�MC�&Ƥ,�&�fh���x�_iqF��z�m���Cꉑ�ƒu���)�ϰn��9�abq$9�in��Z$#[��nGcи��ӈ�7d����ͭ���������~h= ��N{��4,_���@w�qX�M���)��oc���o��-����t��#�ֺs�-`�[M4��9J_������P���6�S�&����)��(X����1l�Aӯ�,���N̺5�\k�b����{��=W�I(��0m��J�u��&�.e�4"Pj����zRnN����ܬ���Ղv�4�������z}QNRT����4�␮�&�c��L0��^��.�̔h�G�j�R"�+��\R��ZD�(���Oa��^��NTŘ�x�].)�p?˜�,'B��SD�����L���>�趽��������R�^$DzKA&����@�B�-[ q4h�)]�<{�nf]��$���C���_����.� $�g�ɞ8?a�[�&���{�b\�yH4���\��H��`\�sS���9�:b��#�M����J�����C�ؕ%��L���ֳ�:�)e� +	dvbc%�G�NI�W�u��P�b��zCB�
�l��yC6ρ'��� �F���x��0�[��@�������d�Q,߻Ł�+�|	9�2k�וU	���ʲ W�M�Eٕk��e:"�/_`��B0�v���T��?|�㘋@|r��#�U�If?���]usi�*�nF�C�m2��B��bAaۻ��8�%�:C~]�i�v������i�ؕ�(]0N`��K�Y��&rK�%���v+6� �j�j<�V��?!,	�Y�Q�_��s���È�'Rp
�	>,�X7�
|�k�"���F�m�@����P�Ԩ�z���Y[h�wڌ���/'.IҤ��x짻T�Qӌ�Z�U�8�ՎT	t{賏Z�Я���= Lh��+�Y!o4�Ҷ6�����٨)� �X�g���'�!� q����u\!�H���Z�� ���^6�� c�(��wɃu[��Q��8�����W *N�`Ck2�����>ȉ�_�}���ֹ,wq-D�P_k�K��Ȍ���V ��@z�اtɯ9Æǔ��bl��8�ypf����D�����'B#��K1OY�2��'���>��o�p�]kÑ�dv�n
E��H%��v�QkԖ��|I���B�m�ǂD�t�����D�g&�/.6�7`IE��?�f7�2BJ1u{�
��$�g-�8U��֮���d ��,8�b�I�'i�Eh�/�>�����]?�pw1=-9��D�_:��FGi�@q"S[ȹ� �3a��tkf	ߍ��@�����42��%:�̄�u���RWH�`� ��ԭ �W�����z�A���;U�Ϊ�N�G6�j���U\�1��>n��X)��f�����a�g��w7de��;CY�a���o����=��G4��f'agp��k"5�6f�G8^��:Ȝ�u=�?��F4�7ԗ[c&:g�5|�q�Q�[�/2AD�;n�������RiV �Gb�f~S������/����VtI��A[���n�r�\
h�����-���HH͹+BDz�z��t+�P���U�Q<�YB�h��r� ��t�R<�&�o��+���W�������?���Z��N����M���{��.#�wt��
��b�� ?�8������n䎼�0F�͵���H��[��&F!�H3�Cm�s|����!�C͙�r� �9��?<5(l������3l�F�y��^���������rU�
��'+")އ��cRa�_�?Q���G�aʇ�4��yx�՚�	�_�I���F�1�E5+L��X�?�g$��ov�m�"��6@*���"#=�ڗ=�Y(�m��5E_^� hC{ԑ���0ip ���t�S���?�f1Ɨ-�������w�i�хH�|ޥ?��t2G�sj��Ӑ�h�Q�f8=���JS����v��O�7B�w�/OEn�lh�����p' ���L�(6�IĿ���<�YȮ�IT�d�ξ���2[y��b6U�� 79��WWp�?G��5�� ���}M���]��-L��[�����3�M{'����i�~K"Ld��M��5oR�bAi!�ڗ�8�=?�3~ �|։!#� A�<g��w|�머
��נ���$i+�`+Џ�`Xg��H�$d0kܤ9��~w^���(������ٮ0�J���/&�r������r�K��+[h�l�~�6��~��S�3|�+��QB���bYMs5��� �δ�F��1�~�IR	���h �>5�gAn�?�P9��/E'D�V����E.2��TOXH�s�&���?;s�>4��Z�!�w�	�Im�2*�ߓmiC5�o���n{� �|�Iw�k�	�r���\�0������`�}$������N��8>�	%*��d��wUp\���u	I@�r>��p���q��'�p������]@���m�#�7	$@3��z#,�cF��h�������ҖD�r���h�8, �,۩��'U�l�|tT�s�����h�sf{�%��rѤ�����h�V�$N��b@��{ _��y��mPϞK�B�x�������kK�ŧ^��*����� �9sJǃO��dP�A8���ԊXE&.8�#��a�j��V�iA���^
%n�OE�2ک]"�2PD"�K��TLd�@J���t�����a�q���\v�� �����\sh0����f]�,�!�怫�]�9^4����
C9�����a+$��җ�TQ��X������0Y�gn³=��vPP,!"�~�\�*�a]޹O)M��;��VEˋf^x�9%</ݺ�@;Y�M�1���>!���}�k��1��߉đ��A&|��N!#��W��Q/eؑ�@�\��8����Όh�[����B#��y9��5���Z3�A�a��=���9)�q0��fu807��s��>[�K/�ν����"�k���C�U�� ��R�x����a	����!����C���(���n9o,��i��!����$����q$���_�$[3ڠsq�ƹy7�qN����h���� ��R����Z���/E��|1�4�g��
���K�2�L{�A0v�7D�,.?^�Qc&Zƌ�����ӱ �}�MQ�Q}���V(�>�dKfJi��f�$����4�7���^��Z��Ls,����0��ʝ����G��"K�!�ڋ��m�z�x�=����������U=bO�A��Ċ(�.�VD�Xq�c�ēY��%[)L�Y�Ɓ�I��v���sm�Z�J��h��]<�R�qa �*כ�U����2����d[��cfQj���Y�I�==�y�1̧�p�#�<}!�	�؂6�#���plF���
�p�D�Ѻ������%yw�����Ly�@��_RJ_!*h@m������r�?N��%ݒC�0n���g"=��x��3����Yc:��y���s�f��I,�;g�w�MK6�e�LV&�"��O_pm 5X�!l��I��h�=̒O�t�K$�,��T�v��	�T�_/��nnY^͔EI�q�����͐E�wܵU}�f��2��7�MN�`�����l���5R@�;d���{#�#�N��e/TMu

�.��5�2kw�
RQ�&>0&l�e��fJ�%���Z�Xs��bt\��~v�Z\� �ޱ���k�]�����O�z��5��c�A;�]OiK�_�����@�kK�:=�d���UlrxBHl�|���O8*MJi�t#T�_�6�����H$�Y��3��H����B)�_��Ď��hlw�<L.LT.��57�v�Y�-�I2w�������y\L��8��N��o�'2FM?j�vs~�3F���>�ڢ.��J�&	O�]��C���]�M/T.S�]l�ձ�Pp��L�aL����`��)8��f:it��<SqR��d)!�n?�m�yN���#�xx~�]��;��l�v����%��RMpH"(��Q�ǧ�Y�]���f�2��P	mņ˗�:Iu�D.	 p� ��k�#W���+Y4cw�Iʗ^C����I}y��&N%�����P�D?5���"�İ 9�JŗC�P��h6&0nPK4T'x�F�Q��I�5X�&�1m�`8X�ߵ�$7@��v9��O�pJ��=2���	+�^����l:f���G
I�:�����x�H��t�KQ-�g�x�{ّ���n���g2w6�t?|�e�
0Qöo	��VC1��`+�b�b�"d�6���-���!1����ӀZ�������(>�t�	�}���x<y<�&�uַ��+��o��ܕ�[d�2�&��>i9� �c�}D�Sa7���ORR���B\��v�~�>6̓R���`��jܐw��C�u����4�FB7߽[w�R��$�b��{�w� ��l4+����1��.�o溞�I�P�bOyT�YS��m`��(��2*E��!��b��v�քT?�(��U��b���%�գ��&���3Ex�N����L�fմ��05���;�XQHX!Z�k7+�mV��|���k��+9�d�:��iX�%:�E2S�!?Eiz��bb6��K����[v�K�7��P<��&�90�LMf��(��'�daBIc��/�6��f�y2m�}�fÂ��ƚ�1�H|��O�+:��w��ĵ����c��`@�U�o�%����K�3k٪j�I�֑��XPn"}�X'�R�L��P*�� ��~1+d*���װuO�7�qR�A�_\��}N�#�5�-��_�HY�VX�N)q��g�����9n�+)�hc����lյ���$3$Gmt�n`��a sL�>H�H�yu�8~l������&*;�>~ā��m�a,��_z�Vm$BV_ ��GZ��`k����.�?�d�r}�^p&"RD�3%�^�ĒZ������y��wаJ�Q�w�vb%s�֎��.P�Culv!�_ָ�ob�,y�,m���[��0���n� ��s�7�b�3�,s��?�\�]�)�
��өINUm��'Z=�ϩ��xRz�N�Я��7��e5~��\�5��B�b[f�����5޴v����,��_δY��bVR�q��l�9�2����� .�[w{�
���9^�HED�m*~�_P�H/�e�x�`�D~�����q.��.���xw�� ���	����!.���
kD2"��Q�As`%ҷ�E��ʧ=�E*���-c��!A�gL�RLѸ�,TH� ��������yX+��a,f��]�Q7��4_.�����gf4%���R��Bڎe+�%��'���@f|��Hb��*�<�F 
ɩ��*0���tgeeAfKH�s�pL:���mI�ZS# �(�X?�B�
���臁[���%�+[�Zɴ)-5�Aw�h:��-&���p[CC���_�IV�M���(Y|�90��o �d�%��.l��@|RX�{�C��Rp}� K��QU,����03��j`K'���y��\hI����Ò�z�����1;�tst򔰠 �^�Ѧ�4%�"�jRte��n�b�9���j���n����g�eQd:Y�s�h�I��������a�P��<��2XN�:ɗ�,Ea�� �y*tn�~h__}�W4bEH����;I"Qd��TJ$��	�� x�Q�t�#̤�>&��]�o��O��j=�k$N�y1��z�5ٵCv��w���!�|��|�0�kQ��:�m`��,.�s�d�l��x�Bτ͉�}�H��3�=�S�e�Y��s��A����[�",������1_�P�B��">�"���i}�\և�M�5:pq�JX�	/1��ޓ����N�/�n]>��ؐL����_X��V�/0��-<�k5y�L�Gê���j���cM�j����J���(Z�!��
f"��7��^@�*����������:�PU������ڊ��IO)E2����,�&t59��~����F���P'*#���G�[nen@�⨭�'y��T�$�,V����&��ST���0�N��bKd���*�ǰ����n�3���ߗ����H�������P92�'BG�$���$'�V�;���g���p;�!�Io.M�zC�r:��
=����&���_	Jx�Ɋ̠9=l�ᚏ"�u	`;��+���]�� _C��:S1��t̆$isr.�?��m�3e�n	ø��D7+'C�Ob*T�yR�绻���t�_���,f$g��˅�
aҪs��҂�h�R���{����a.��a�$X������'�)	�2�u�O#+]�y�`���w���^E����� wA)ܻ=T��H����J	��̦}���;�t���ͤ.�1��0�%\1����_�owe�p̐��PM1=�w���,�9�����*Qf�.�Ob&gi�7ύ�J�3��Y��a��*z���6!k��ʕՂY*����3V]d!{�	iQ�r�{�_0��'�4S	&y�)�2��� �Â�Z-scZ��$e�6_(��#��6R��qf�f�,�� ѡ��#���&�S"�=�s�so.E##�)��n��r�8+9���Tx%{�����ꤿMUU��O��C�3پ����0� ���WpI(����t�@���E�D��#��k�Ln�8m¡��	�S�N/�#n؟�n0�jߜ�.�X�珺"�!9���IzE8s��Q�޽F�ݴz>0��͵�I��L�(�QW���W�
t����e��S����*��-kH՛�$TQP�T"P0�������o5�><Y8��M���]90��d�_;�F�R[��i�,�;	g�ݜ��ф�P^��2 ��_l�����#dEEsa�g�-8}�Noi��D�t&MJs#Ƨ�+{e��a�jgO���!�3}W1Fх?[3;�O��v
]6����}�|�H��&�*�_?�i)L$����6	+e�s��&
�c�l�>	�;*f���*�Y(��M�x׋5��r�b/�z���;+��9K!s���*~�;�ةx����. �؟R��h[��J#	%:c�Dw/�������3�ң�x2J�'Vg�7AgN6�s}+��)�ZOg���H�$���U�K���Ϧ
������7����pl{�1y��'zn�c�^Yvy*&��=ݘ�6xsf@:d����x�Wr
2%�6��e_d`k�N��'[	MG��!��ak�AqPf�w��B+w�I��@����Mq�i�՗]3�|�E�0L����޷p;���CV+�*�4�z����w�膭�7��wj_��ʸXKO'Drb��?�T���gU�d���u�Mh�3%~Wx�*��
�Z�Tb�84��%��T�1��a��鹼c?T�����c�����ch���n��lg�B�rР�F���Q"�n��qjhk>a������fi�����N�Y����#	OͮNpP��5������z�F�m�נx��k�JU�;��9�&�N�}�v��!�il���H4p��h�����G�BSkȳ*�ll!���2�KU�}0�#���Ac�<[���&��?���{�������G�'���w+�T��[C���2d�Dv�ωv��� S�<���I��N�.g _��I�˱DK*"��*�P9�w���n�)^J�H4�q���֚
�׌t����M�u����Y� wy}� 0�J�����'��\ ~ �4fWojT_[U�R8{��$�H.f�$��5i��_���0�h���ԵMhJRU�Զ���Wʂv�-	P�c�h���4�VO�UTou�̲v9��}�2ZZ�q�7.d���]X�����2�K�L�n*�g�	Ƶ���]RcT�#����xȱ�)��q�y'�Dk붠b���l�W�gtR�����\ePReӝ)PVV9�طY��@`ݪ`\�&8�>�oP��`���%��Q�9,�R��vؑ�d�ݓ������;�h�#��1t15���,�}�K�ζ�>FE����nL�s�RJ}q	�����;�r�`�s4���V��¿�M�b�x��������YQǌ�m����#���fZ]Ӿ ���=8��.Ҷ%#1\�zBo��N��Ft�<#�9���WJ�%m�T*�:��*!;���O~�Xw��nյVw����3V jOЄ���$����3���=�[Z�<���qZ��m��9����|�g䰍s�S])l��=���D�ƈ �Q(�T<2�\�Sk�7n��h�6���
�#}A�
��\2�E�j�ECaX0L�&���.8����,��'C	ʏ�D����?4�,[����q�˨3a,��b�j��,Z^e���l	�{�_8�m��Ao�t4رE�Il�����_J�6njоv�0)L+�[��!c`��7z���\����bY�tUR2���r���o�)���F�`Љ��:3�s ������B�ʏ�d���V4��n�����fQ?���:�a�,J	3LЁ��e���!�_�I�V���+�Yg"����r��/�:�7f�Yr�55�R���=k���1<�)�R\��#Ʀ���W����#oXQ��]�%�����h/nYY������T������*.̛*S_�����#��L�[�ѿ��У��6$�=^}1!D)]�1���p�*���*��׃s��+=�`��R�4B���Y_�y�
-Y�Q��;Pa�&�@ '�� �n�L�#o?�0bW"�DTV�3����K�J�ޕ��-�d��Y�v��o�Pi
�靆o��nZkl͘�ԅ�䶔9�\� \���y��Ƥ���V�u��є��G�%z7�����o��xb�XO�O��Iu���
e��m�=���y����'>w�Qr�y`�͂�����(����(���B	$��e��@xO�O,�#�j�(� '�%#t�)�'�QH����m!	��M\���$ή�(,"��ܳ�:0Oe�q^9զI� �x��E
Oh�2tn��?�-p��ll�Iu
�\ߤ�^�%�����ǽ�$C�'�d�j�p��y��?T�*�����HB���ogN<k�gL� ]��s�v��@?\� �d��{�5��HC���6���0pT�^���t��71� ���΃��L$����)K�l`�NLd 
껤)�ڸ'eFЇ<)��Iy�V��+(C�6����ݩ
�sS��G�QӊM���
��`��	X/	b��&p��PW��@�P�s�N]�*~���9��|w��<C�ݘ�p�~� ���4˝0�	
7��4��h�^ּ@ϝs��rdT]�ɫgA����!�F*��3���:�{�OQ�r�7�ZF5�,�z��B�q�?��>��Za� ��zجp��}�ى�v�c� �Yan�&k��l��&%8���S_f��]5pP׷�ex���`e�Ok#�����'�>�K�� ����e�ũlT�����#_�3ef<�ʊ�<����%V|~���&��8|b�Q�&�`Gk����O�7�↔۶��'O����𿳷jJ�����M��*��i�;x��'�4�ɚ����q�FGS������3�&}�M�Fnz,j�r1�<_��S�r���,\8x��_5o��h@�c��]��+�Ɗ-)�3��%�J�W�q�=��o7���R�wr��T�Z)|���r:W	�R���^,�<�-�ޫ�E7�C�f�P�SV���,�'�3K!Lg�"���+,7��A֚�fsQ��Nz�&��A�d�E	��P�#盰�r��x�l0g_�^ʕ%�:��P�u����.�p�)��M۽E��2a�I���4f�ێ;6�
.�xW�ҏV`K���z�_�����b�)+T|�|٫�o�g��'�O)�*u9ed��y�C��q���~~J�J��1���c˛�����˺q�1�8�z&E��&j/*���Ӆq!q+�WUK�W}dbx��)�|�q�L�ΰ�ZO.����bc �u/)�����J���������59�r �W:�%-pPׂ�}�ky�y���0���e:�*����|d�qK$/Rh��{a�?�_}`���g��D~�������Z��aB�@�I���L���+�X,aʺP�;�*wthR)Y��\=.J�:)ի�0	ŒЋ�,�`�<F�J�\gE�P�Ā��W
��a�[G��L���������(��<��G$J������y���߷s�����l��6Hu�SK\D��1L�='����� �3]��_7U*bT�Q@��D俘��Mi���&>�u0��|��&e�[jc+{��gNt+l�@�b9�.�as����8C]%y��Xg A�5\D����٫���]"}5���:5#��-�1�"��xH�hn����O��� erOdī��E��VB�	�d�֜�	u���]�V��P��s��a��_',�M	5~A�����L�87(���
}�NP���+�|x&�e£�cBNd5ˆ��.����N��5H+��i�ތS�a��3S~X���&Z^�g�?���&��qhG�$!enU�Db|��WE%�䍧�@����>��wJ����]	*�Z��=ٝ�R:��,-���$ {t����;%��#z���v
��a���'��VI��^4�Y�.����]�؈x�z�S=f�vHj{,�*g����a�	��ŗ��'�����.�R#QXk�D*u,�};��&��4U�	ʌ�I���?e�ڽJs���Q��bc5+���Z>�޿�hd#��|<���������9�/���~_9�n�|�q�K�k���e}#��P!*8G�(k/�.I�����ik�c��p��*$Bk�)6OFg���Z��@tl��k����'�vJ!�(&$��0��7j-e�?pZ��f���{,&��
�mT�gDK��3r�&@��T��{(z��oi)t��U��h�$��s�I���NJL):cM��[R�G������V�(ri��d���RP���/�ty�bܶ-�����i��!�K_^���ɽ�����H����?�vkD�9��� c��\��,6t����3�>U{�d���[�������*���&=u� Y^ck�c�	"�-@�Y��ݤ��-�'s U������`}_��������g����bl����=�z[�Z�ȵ��OS*:f��ܫ-n��b�����? �˻���ޅ�,�$�0���@E�5N
�ظ�ӕ��-�l�~ܿ�個C�����-(R�y�(�A��7B ��/��������q�,K��0�*sѬ����B��@�n�����\��B������%��mݤ��iN
x����Z��4��\��~�����h�+U��iﺚ&c��&e�inX= ��b+�ƀ�=�9<IU������W ���;�v���d4��֧��Wj�z��ɔ/�r_`I�v~w4�HJ�x�[��g�Sr���;!E�,��Q�}.P��q_Kͥ$��g)��ӗ�gu�pdXN҆�����X ���Q܆��?ȇp�����J��`�V��_��M}P�����vb�BJ�e��Z��09��F��
đ��*�b�&�����H
�Jm���"u��ء�J��F���˗�`b{E��5��ɰ0������&��<�bU���e�Y�
��`�2$YG�,@b�l�?0����h9480����ONz�h��Mq1�J}X{��rU�ËU�βncL4Fu��`�&��=W��(0���M��r�݂q��Ԣն�bsE�"�3Rm�\�X��HC���I&
�ǭw�x�,tƎn� se�PL��S��GJ�5Z��79xb`�_z��j�oj�Gl7:�A�������[�/�J�S�Vg���������%��q6�d�"�0�����Ȇ�R)�# ��{q��������(4h 5�O��FLI��r��)V���x����w��5���(�8���2�0�Q�"w�^�f�P;9Z"�.~<p�t�պ�����%}���[AN��)�t2�O"ʇ�Y� EB�iìa�O{���?1�pf�������âb
�z���;֨���ȥ_�r.�!����&�^5��Q�RhE������5H��Za�١�OC�5���uߘc�]ʠ��z����L�R�8������E�~j%������	�iL1.�d�@�H�����f���M��|�����8F3�k {f���đk̜2ξ��� �:X&��kM��'��-ѯ����݈|p�mv�%�/C�4��}��!�f��
�-m�1=fvũd�V>p�pM[}B���o+��"XJ�x�,�Xq�B��gaE,�1��וJfdxG�J+n%o�be�d�$�����"�.��L��^+� �i#E{�����e��
|�i#BFd_�V�D��h�.��[�|����;��~o��o�Q�r��惒�^��ڇ_�o��v��0өU�[�����W����|�eeD�_�j\��%I�Օ�ށ.���գK}�W/,�*���< �{���(��֡?;��d.�N�M�D',�7H�)�y�Tuz�eLʌ��	%�T:
��Om�ޔ�wu���鞆�z�Jɴ����0������=y����
z�";�]���B4b��j���̀��c��&�WCM�����#gv�6I�j��m.��?+Z�g�GY�Q���W�<�_�ͽD�?��BA����zTy<����{�\������x����|��/���wz#$���,_3��r/"k�U՘�F��֥;��4�J��[�_���ׄ��U���{���-�*
x�b�Z8�G���%�<�8����� C'Z}�!�`�]�&c��Op�����8�����]n�|��
��������A��Ke�鎳��mL�h��*+J2�����j���7�y�K�a�Q+�ZP?���.����d�����Z=3�'�lQ^�k�H������~t0d���( �V��A����ʆ�f3׌ =�+��fX�(� ��a��/f%8�J��.�քt�GQ�����`����:S蟥n���;��%�Cf�ТW=8�i���X�:��U�S�����;�+-L��MU^�DDO~m���f4,nýt�8�"�F]Է��Ҥ������z��bY\��'^��۴N�~����A:]?? w�u���J�m+x#-��qN�E�3�%���cc�vv˦�o�4��6�M��L����i�81�kP����h$�Su�E���J2ڦ[�Q�~1*�/$��B�~�P|�l&:cQu*��ڽx�<ҿԚ18�UG�3A��0Q�^U���%T�2���{
�j��;m��@C�,e���C�3�B�-.�Ǚi�z�N�'8��4�W�׾�G;�����/�/2gw=���z"��4I��Pǽ�B��w��4�>9F%��,ߘ� ѷ#;���[���g[����6���ź
���i^�x gȮJT��v+Gѹ�kzv�� �����41~Q惴�G�l�<�X��9��պP4B��cݮ�<p2��e"AYx��7�{d��Z3�hu��EK�4<�z}����V>���͘��u��!#�t������g�V�,�u�5r&�r|N�\8�R��6�������5*�P��!:��iyw_�%���}��t��4G5�i-Jqg�{��OFEh%Ȋ�d�j���9I��F'�4��M5�{�'X2ǋe'c�5N�K�u���jo�n�C���>������k@~+���/���n���������EF:6�-g�(p#<�G�C�����"�@��yڣX�?�T��Z/O�̖]-�A��0į٫<�(��{���t���rFHۍ ]��y�(*�*���D0�I�E�
��=$c�&��T�z�0���%�SX���n�์)��PBD[���g�y[	�v�v6�*��52����������=Y��vZ�f��fE4}B����'�9��a+3=�T��T��G0<����H�џ}�Q:D`�����_�ߢ�~���>����0bc��bb��Q1�8�s@ᙽB���):f�c�)���]���Wኄ:��M>��$��D�rW�m0f�DB�C��C�Uɢؗ�Z#�l{U���[��Rpl��,���L���#�YL���a3�����L�G��;�P,=4�E����p�~U�(�Iq����s��P/�� �NF��E��q�/�2�����Ov���\��:�<W���w[������TYkw���5�j�I�S���aR��b��i�≻7�`����TZ�]���@��DS:lN� �������,X�ux'��1��f�HA�9w@7��6�����e��jq���s�.5Hv��ߴ]ޞ�Bma+�j�*!p`?��W��پ��@E[������l�o*�%�LIY{�vJ*�L����P״�wv��S�@���}���Ad"%��!�E�P^K��k?��8�d��y�z��I��+kGdnZ!�"'��~������d�����Ne��C�8uPH$"ޢY'>E�gP3�n�#�9�C��	[Ç�y��9� �Ѩ��v�������7������O�?*dc�J��*����L�GV@�}�_f� �'��Ch_���0�l��<R����L���"�����?g����HKtT�`Xi�s>ԑæ�Y'�^'�y�h17yw�jhe5��:#��$}0Yy-Y׽��|��W���0{<��|��ﶳI���P��C%碫9Z=4f�T�8S��P3��q �2�!,�{����c��@A�0b�B߬ɘ5�4%�Ȅ�-]X��ƂA[�G-�,7!BUs״�9]���p��y$%�6��*��wmک���D�9�A2��PN� �Q|�D�$�}u�L��@Utվ�ф��O�5�y��?�FG�J����X����^�*6�?r{���'��01�K���T{�&�j�d���������w�Q�S�(�о�����::��JꝤ>4�7SʓD�ߢ\�Y\8�2ho$�l(i��������41ʃuy��C]��i>y�g��I�c���f�uQ!�ל��z�Ty��?,t(��������[[iiL�G@�3]� uf����~;d�c��ɮ�����3q��f]�W�#��'�7y?�f�"���z�ұ뫼�&@�����.	���nI,1���g���E�"�)L�̋���~qz���4��!,��9��O{�[*�am6���.��W'֗�P�S/��s"J�	�a�o�Vk��r��#�Y��M�M�ً�7n蟒�b��?=>	2d��k��`�!��~:��;Sv��w�ݣ�i�ь��5c�f8�(�y�n�����U�v���Ti�O����j���A/���R˹YXl\�9��!3w��wL�{~�1�;D��:�h�qC&j�a�#,B�
����O:kC��:�H+�wm�W��(���>�
��c4�<��HF#�!�nV�r8z�g\���bP%vN��Y����+��[z�s�����l����z�����)2�ԡ���X{�7��A�v���^��1�wdb�i>�}���X�YQ�5C�#$�c�4�8@��p�w�gY囉��[��xn��n�����ǲ�[�L�H�!����ս_K���!JL^�h ���!zn�wX��]�c�XP��[��!$*%Y����G�����װ�{��Z�

��<��g	 Sx�_+��k*�٪�lAi4U�2lTS~|qĔ���W�ޕt7�AQ7W�dQR,V"<�vt�����Q0�nEҼ�'~�?(��R?k�:޴�Q�"˟z6�E���hPڂk��}CɏV��@� j������;W)Qf��yh{f�}^�h�<��a$U�ƭke23b�^_3h,���7I���m�>$&�ݧ^@�84��2� ��P�d�9��5������+���8U�;_5qɲj!������*�4�f�K�5���H���S��Z+�} �҄���C������o|�87���O���
Yvg&΂^28���T�<ȩ|e��ܲ�M��V���l��:!������:STsE�&A�s(�M��KV�R�vb�r(�/d���5����G�U9�?�=�?i*y�id�S��{s�/�.�;'��lG�U��R[u3�
�DDV�-DDR�Աx���eWkrW��)I0�c뜵a�R�V���_�u��R}r{�Ɠ�6�'���m`�.�c�@aLѓ�(-zˎ(�Uz&�;����/��d�n#�.�H:��6�[.Ռ<�HD��{G��� ^���9#*�wQϰ ^I�{�BF�\k�DUf�}ce�(v�s^��,�M�)�O��X�Q�^�L��K�,c�fI�t,i$m�KS��. u� O�~BI�Uu,��\��X�X1D��#�!�a&�9�Jp��*xVp��
z�9�JB��Re_�Lc"��FC���*�[�e��'$y
ϝ�h���-%�9���(����������Y�Y�
z��R[��=���o��L�8�$�z��3P��x�z��Ti���J�=��d|�:�D�#�N�587n#p��jI����)%��$�H+�ӟ�j�Zf/Po�&ɉ�"	vi[Fj�c=PU)LRX�AS��=CQG�t8U��t�Q���k�ڠf��*M����3�s�O�A׮o����i���3�i��f�U��&0��[g�54�V������NH\���L��9�q��-˚��x!�gl���t)U��`��D�'�#w��m���M�yQ�&�3Z� �� ���0�0rB�5�z�9g+�����/�#����(�G�W�z���
�&�c�v�[�ߡ4��oA:[j��`��`v�J=E��--�7%YL�n��d��⟣�Z��)���$-%f��p������� �!����`b������������L��2<YM�{/�S[�QBVSe��7���������y�?���Ҙ�hl{zk�0p��@\?��xZ5$S,+m���CTb엢�{�bF�ȗ��y�����R�~OF<a��d5�	�����9.�3�0���c%9����J��u&��0d����ڳ�"�S<��	�=g�-��j-2y��hY���(���';�Ӹ.��b�+��Q��`/ָڙ�`���ԙ늪���=��1x�L<|�LN�k��8G�gI&tP��l�Cܺ�%���p�x��*��Hf��R�����h�m�Y��Z�>��Hk���`ĳ���R��w|/��'�	�-�ap���C$�`�/��A����;O��)[��m{Bx�T �E����dI�`�C��B�v�М�p3H���F�$J��@���X��I���@�pjS$B��;fѦX�@ǮP����m��K=WI�P���+��!����{���U�8+���R��<7���7�j/o���'���-`��n�[�����5z���]x=5���)�e���7���4 ��!T��Ͱ�bkҍ��ݹ5TCC{�}�e���i���A9��RL���)p��o&y~ξ��� :�~��d��og���%�5q^�󥃩��q�����]��Uo�N��h:����Z�t��k&y!rHY��\c� �z�C��i�[Y��@i�admE�[��x� �M��d���z_kc�&sh����F�z�V8����˭��'t��Qh����(���K��{�[�5E���8��J�K��Ȉ�&%�`��r.�gp��d�nb��E`��7(��[����>"y��י��������xr@�.%+�TI� Q����QRxB����{[���Ŋq ��hS���K/	����>�kR�g��-$�OqQ�PL.�m�? ������M�>)�@)A�����4���xƿ��jC��9sA,4p��ҦԚ<���ʖ�O�ߓ_p��J(�k�	a��Ϩ|�K|���u/KE��DO�T�##Aal}_G�Ib.�*��#�tq�E�7�=�y�=欃��Tǧ�ǘf�/�.Y��i3�6�q,^�_����S�B�
�פ��9��Rm�B,_ӿ�z]�v�v$�!�e���ic����$�@�:��I�NX�8��l]P)�C�B2ڰ�X"�rg5�A��Q�t6�0?l^9:��������T�JC[uAI��� �����HȄ��e��G��V��dlD��{�m��ir:R��i�%ík٢*F�;�^��3 �g��9o;������a.�N���$�U���?DG�ݭ@��X�<<�^ڏ�"�QL3�E�h@����!�sή���1t�[cV��]B�����^C�~{N��k�-���VK�SNB�p<9D��L;�ߒ����y,֩	�sU�	4,�m��4Fc�Y�H�=h�X�d+�gB��F;X{��~�z$|��ƒ�I��J�]/!��g�%��D5�UQa�Q���m���+���Y�w�I5�8	�N�D3�W�'8�7-v��o���szE}��g12�Q�n��,DrT^��U��o-�k��mm~��3�k1�ӧp�\}H��G��-�_���i�Ֆt��Q�@�P�B�
%jr�>��� �:;�m혶�l�H��|���C߾�2���Fν���%�Z���AL�4��.�,���PXoF�b*
�(Q��d	�������8�h�j�>�T܈.o>E޳\���X2<@p��2<Q2�Q���C<ll[���oA�|���K!���� ��k~s�Mm��[�Zc���+�V*!�1�������_Cfi�����6����]j	&���`nӿdS��s��[�n�9H�����k7�΂\��U�@�T�v5��`�'�N�P�|N%����~��x���wM)J_ҿm�y6�,�3���ke�.5ş �]&��eW�Z�tU���'�H�QP�yOp<�p!��g��[��I�$s���1�=��T�"��vD@,�EP/�m�.�|��~�h)0���6ǀ�~�0���<q悳��աDqʾ� b��"�ԗNOĮӿ?-��cF���n�ol�֨�m��P�Ɉ��S�~��{cXŎQT}�
�����L�m�mۚy��S��3��&�0��]}�3g��7'�?1Ÿ��J�t��b���ܤ�x���� �F�"��ȜU_�����h�fEh�n�6�ψ׃U�^��~�!�����X,��syJ�:H*ų~�i�MFq�M�q��m��*����}�veD�A����e�+͛y*N��u-����[�n��ul	���p}��O��M��Cf(�pE�fF[S�\<r�T:�>}���]8	��J�^��`�Gj�r�G�0�ú�7L��q��u��Ѳk��+�ěp ��a���:74���9M#a�eI֦��S��E������2�����y�i��r
#!Jbe�!�:�Ĉ*��Y�{|r�Fim�Ջl60a�o3��(`u<�9Ht�m��0Ŝ�?�<KC��X7�������g�pWz<��<|�r�T��U���vY�l�r5��q F���C�}p*�GA��ݷ�4����)U}�ދ ��꒐2�Sf��G֧鱑v�y5�N'�s�2�7�^��:y��=�+�kkz����M��7��åP�V�5��(B��Β�����S���p]�[��F���m�(w:��$�l1������D���H�f"�2bS��qO�|D>P�]���r���{G���������`��Q,����i�gIi&�FW[k��肽�P�n��xeơH����7Ar� �\�Of~���� 4��^=A���!_Y��
�*�AN�;��g�뜽�xX��D*,*����X4�S5
$�-y��+�A�;Lo��}�M{�����ψ�b�I��M����ɍg��@���(�X`��?�ޤ�̱4��ӌ���խ�j�O���o���Y|��{���9�$������ ���ݦ�hD��,N����Z��w,��T*�2��Y�	hy2i��2ꥍ��^S
�7_��\O��P)�1���x��;�bo��L'�0b
QKՊ��->Ft�~e��M��l��;Y�\g�@waj+��/��epk'M�d�ˍy��*���<���-]��Q�N3�x��	�!����rV�C<����7��/���+�n� |��>_�(��S"���P$:]���E��f�m�Xc��v�C2C��1r��D�������<.܇�2��(\A�{/�?�,��؆�g���f�b5qaa�'�Y������ԜM�G��$����tݴffO_�뀳�1ei���'Þ+��*v�x-ݙ��5�:$n7Gٳ�*fKd�{�e1��K1���	z�����^y��C�,��s �9�Y����u�ZzX&��B�c�ަ��E5���:a�y�b^�|㰞�GP6�2B�"�i����EOc��a~[X�-�5WZx��?5
���UU�����ʟQ�g�2��7M!��.��X���(>�a���gʝ�廠@8	�]\�U��R�~Y�s��f-��*&������ln
~O�ު	��Օ�4FE^�t�y�<Mt�$�,X���fA���9��d��Ҋ��4�Bu��\������7ي/�ZrO��mG��R�F��[���}F
�'l�����O��$]+�a%FD��7���Iu�c2k���bj�%(W��(�5�!��*	ěsx	��zs@��i�����jjQ1$y� �8�g��� ��Iq~Qehͦ�5��+I-S�����X�@
 ^m�0����I;�"B���6���x8.��)m��E�W#�w����f��C�3T�=�4ն��[e4������-'������+�t�D�#��cQ��wKV�Df�\ȸ���MƋ�!H^��bȔ`C\y��'�q<��#|Q[��}i��EԐ�r|��*q�3���g�r@�������Zɝ+ �}[<�c�����v�	[�����㽞 q�˱QH�N��w*!��X�Yf���2;װ���M+�<�= �߁Xd��x1u27����Ѥ�,mq�>>}������u%�p]��P�몣�&�)Z���^KO���D6|����i�p��B��ɕ��^��ې^��)��4:�t�&Bb��u_u�e����`�~���v!�|ޖ2m7?�ڶJ��`�,�]ս�&y�,�t��}�I3c���
7�{wd�u0�ڴVk��V.�� ����A�2$���T)�%�_R,x��I�Qb�8a��A�o�Q���q��פ^�����Um���p�[��>AS�7�T}7�[���P����P�R�|d洅FQ�)(4@(�8t˹sw8M��i<*�!�X�:�0Pt�>��¿�r��l����C���h���uI�IJ������\�չ���������`~.�Ji�t������,�&�=������Go�R7�(����]1&΁ӷ�?-�&��!��c�dX��nFd��;���6� "�C*(��t�d�H|��`#44�	��d���l�#�uR�b:9�'@���@��]������%9�(�#R�ۂ�^繆�c�4	�k*ՙ,����'H�ү��"~k�3~����d3C��׏ä\V�F.��k"��j��_ �"�̝'�'U�E�Flwc��~!�r����1���mT���v`�_�	�	9��-䏸�(�V�bn��A�t��p�5έ���dUQ��ig��V���
e}iTS�E~�BOO���0�����%�F|�J���J>��'��$�2��ҨBjH�fﾡ�:r�i5C�8M��2���[%���`��=L�Oe�"����8�y����f��'��<����P�0$���А�)��1PQ@J��Fe\�^�0�Р�x�H�B����.(�(�y$�G��d�Lj���,Ma��Sf��������p�aY��zb�V�� �P�LJ��dU���y���T��W���WZ�_��}쏛�H�||�'�+XaTVxk\��(ܓ��Ae���������#�
^�J&>�ߓ�͍��-܆�(��dQr���_����$���#K����>����խ-q��/X������2�ˉS�WB�L�r���?z���7��8����.R�̵ּ�o�ä�h9�����/�P�r��>��1d���8��)2	|���d����g�ȱ����8��'��ޘ���#�0]��뛸ݓfbƖ�T�]�F���l�W[�B�*�0����L��刬�Ulʱ�]K�\DH$og7n$O���t��O�ڲWrf4}@�D�^��sC��_"���.�ƖN���-�4�� s���4ŧ4p�%|t	�=Y�,]BQ����Q��#�d~E��ۦP�xѦE�|�!�Zѫ�3I1��o�<�_�>��`������!	S�z���8�
A��3I#G�E���q�k���$���G�Q�e�9��.3���Z�e��҈�}�7EJy�����щ;
����,4�+�e���;5nd�:̽�T5�Vg\����g����hpr�NF��O�|1��*m�L��Ϡ;�l�[�nT#on_�w��,�ٹ�P��^//�4�
$�C��9Z|Q�E|ר��7�)��<��'�A�A�1��p��ޣ"�ʍ!9Co-��"�x��X8�?L�S( ���v~�z�{��C��q��J95G�
}�d/�rT^"�d�]�������/��Gq����.Ztd�Xi�D$�d��g8�z��4C�v�P����9�Oс0�M+ l�w�e��5����f���ݔn�+�'[�X�g]�F�-���u}�*�c� Q�y&�[p�LT��>VJ,�<��3�<�������ET�I@�O�΂�\/�8o9�/窿�:K��@�)����|ܔ����cx&�n%�׏���ḙ��^��%iDi��v:?А��4N��c�����(gQ�w���ZՇ��o���:������Z�ExB.��N��M���̈́��*6`������L���R�tTBF!�0�s��"�pqc�K!�-�P�PIh*��m;�~b��7�Xr��Q���~୨--;���������J5�&gk��������(pzo��lC\^�3`��z��(�O��=�"&�y]�~}<�)#Ǖ
���	E�TN%�c���#\"ߔג�46�����ʏ�N�${1��6���(����4�m��}`�;*O�i~6�tV��?��_<yJ��B)Vz/�������"���Ī�ꦛ�i�,`PL�A�O���VV��:��.J�7ꙡ�5}���O؄�������	,��ˮR��B#۾{�Q�#J7���v*/����;nM�+��	�_yl�C��s�ղ��j�yn96�.��ABE����D^z�4O�@��z�Ҟ�����*#L�!�fE/&��`0�5����k?كP���S6:���׺�F�p�Ql9M�{��t8����&��H�����lF7�w�� Aҁf��#*>�F�S��t���҉���tΊ�?W�к����f�a|SP0��E���\��ш�����\/�7���$#l���g����Ợ	�O[jtZ!.3I<�+J���aj��j]�����R��u�h�Ԟ�}�i��'����3��,�����`���6a���D�΋2q��M��P���abŽ��3��2��p�zmU�� M���y�(�����:���}�ppV�Д*�Uդ�U;�~Tl�NԄ���T*5��`9����}|=���Ӫ���f}N�\obQ��N�C�H?:��KW�.8- VO,/��f%:��6���]�J���r��ܤ�n9�|��{:A2��L<z�>��M��ڷ���q�׶��t>B�Q��64hM��6��HOG$��61Lk�����fW%�	�'�>8�-�[/��=Vy��=�tۀ��̀�������L8Gj#���ɥ-��Y֑
� ,�c%݃��{�����O�d��5T�7���&��<S�����|�7:O�q{r�\TbIO���8\-;	7��]h蘳���Vd�>�*�|�N�-DI��Axyı���F
/��.��y�hx~��q����ɲR1�YUR(��M�Fv��c��t���X R]�e���%�#5�����f���C��
��1H�P�V萋("]O�ꆝϞF�E@�_�	㴗f���c>d�R�.1 �#.����v��f��T�����*h�<���[��ܑ�M$��RU��CW�?���Et�����Q��Z��@)q}�1/(~��H�_�u��ں�H�t�6;{�Q��������`��8w������R'�q�T�_��W���ۥniDy������g��v͌Vh�H�Y����>b�;�����ry��
�@��R@v&WINn��4�hf�U��:���kHʸ�Z]'�O㓤�m�m��D����d�i�iR^��џ���_<B����o=<@so�f���+��@g;���Lg�n��>M�5~�c�:�����PB �ʭ{z�f��,�a��$�[?�|v���W�Ϲ��Q����nah�ׂ�1�1���$��T%�9��K��@򋽞��Z`>0^`<kvѳ���j�6�t9A0�"��\u��C%����"q2���4K���읏�[�ӌ�Ԏ�h�Aꊦ��ver��qk����+T.�hV��-���C�4�C���WIױ"��a�)�x��8��Ĥ�L	�zݭ�E��xO�#*n��e������A�[�0�+��;ƺ~�+}-�����eN*�/��?X��� �����J��a�߽]���
tu��Q5�+an���,;�̨Q���oJ$^���f��n�~8�C���\�����у [s� *�� 0�$���B��$��hH���{螡�ϻb��z"���K����>�������O�w=Bި�k+��$o���KV'��'~D���I�D����DO�.g�G9������h=���Խ�����n��ش��q���7jj��{+�|�h�2��6v�K���l��XA����%���+*��VE�l`�J��`��;2����;)C�d�T�y`�����>a�P��#{4bPk�^�@�e�XC@�j7_��c־�D���(�'�PY���^����u$t(J#�����{��Y(�`q��Pg�K�|��\z�y�1�DF�y���WKL�g�t�._��coM��3�Ϳb�gF�sk��Ѥ�"!��:���&���?�����6���R5��OW�H��%��7Х]���������	0��� �
��!|��<ṱw��b����|7��%>|� �VܾFs�����4��,�Q�?
��:ȧ�((�� ����|��ɑ6Gɞ�:g]�7|����^z������wC�nU��Ra���޶��M$�
Q#����ioi�ȍ+��eKs��6<�Q۾�d6���)�4�z"2.�/H]*S���
�ZQGS8tkp(�H(;�y ��V�!�E�9��Zro�E) ()��@N �q�d
>���k;(^�=�C� �1��IԄ�E�}����r��ӑ(OiX������ާңR��m���b��U,���n��O�JlR���1����A�޻�L	|.��ypZo�R�"���>'!W�7�.��פϟ�0�58o(-�r����$��4��U�������fp�9��z�w��k��EX�����@��1b�����ۓX�֒�;*��[��Bę��_��~=a�t�J��Մ��i0^iPH0���(�~G	D��Ug>O}���mmGz��Ǐ�D����|���r"C*4=�7�3�'�y
��f~y��PM�ȃƩ�0��[��t��!�G����Gk ����Q��O��'�Z�4�����Ql�k���M���u�p�^�Fȍ��r4�@���P�>z��i�WT#���ƚ�d�a�xG(�`���8��h:������O���&&���w�QӬ�E<8��Q���lx�+p�u��B�Sk l�<|?o�gZs~����i&��o����=!�8R�|NZ��)�U���aB��isC>�ژH��=�1��J�J؉0M���anr�2R;I��Kv1���4�}�����(J�2�r!���x+��m�Z�ey�S&�
�Q�F~���#Q(?�-�� ����Lߩe��,V�szM/`vݛ��)Аw[_P�>3Xԕ�|:x�6$$2������ �;~t�IgS�|��E}USq/��-U�����0#�~�^zf�;W�w�'�6b��e!'���ի[F+Y�u"�q�����6u;Q�p��~�<�� �v/ q�^o���d0�LȼԹ�8�w��L	YW8H��i���!G�F����NOt
>g:��h����;ѻ�����N ���_��5�N$'߰�Ԕ��8���0Ȅ�|��{� {�߀���
��z&��b�Al-ŽC����}��Θv�R���S�c���-���k�f\of_˓z	=�i��3�lZU�i:I����<��.���I��,����$�-
@g����`yP"^��.����Xm2"�K7���QY�
�[���-C�gR�F#5]�e�C)� O��E|��d�{�h��/>�Y�B*�2��d�-/3��k��&똓?���;0���~���|F���v��u���9�\��م����n��U�y:UIMU�.[,c��4�\��y���h�te?H.�)# ��_�{�y%'��'Y]�K�|s�� N��LWS�g�p�[	��>��.�����L��LǤ�:+Қ��u��:�}�F�f�� ����
ѵX�Ԗ�8�)��g_�2��jx���9񅓰~�C+���fO����8x��^�u\���iE�H;�����U�2_�U�����_�)�C=����7�����6��ݫ1f�>\ѥq�(�E��I�G62��}q��|�:�5'�N?\,�����71T4긋2�n�?�fV�� hk�{�g�$Hܼ�{�I�3"�k�/ᦻ�f��Xv6<���?��5Y���
ZA�?��.�_��K�:�2Z$�qt#��5���u��9�Ԓ����2�=z��@E�k�,�5)�E�̌�@\�	�P78��9�{�����s�#xP�9E�e�O�[=�G�����4ЅK*�K6Mc��~��������hI����4Ї�h�b?~A���\(��%.�["M����5�	�;,����40tXR]l�D���2G�;��C3�������(dt�X�<-GL+��T��z���&oNp<�T�ұ���G(�(���<��H\�m�1���Q�g���V��!D.�<�д��7������	G��m�����O�}��9�|��7k#9��O�Z�|5'��0CE�(�mཥ�9�}N5��&���P7S��8�Tݞ�̻Ud��,H�G(�~��1]�����g���Sc&���/ن�������~�]����NWy�024������j�c��<5v�����J��{H��\u���:�Y5��=X�W�o���]���j�*NH���>���yejN�(q���,<I�'Lj9:�ϟ��3�-w=d�\���
>�:5ϓ_Ȼ锁8H~����n�Ѻ��{ 2��W�ET;!�a��);\�Gy*�p���[�EԯO��=�cJ�O��� I{1� 3��M�n&����o���<\|7m�7�GU�E^/�1�0q�3��!�\(�9&+�Q��`��gY���ִ������ad;i���׈��a�=lPE�;�M6���H�&7���X�c@MT��74�.ޣˆl��-y�v��y`E�-������a�M��*yO������Έ��BӋ��Z�԰���Z}�)/�?GO9	��ïˎeצ%#soHuNiܭ[�l�.���~n���c�w�~tm�( �F�fY�]hi;Ĥ��$����yHn��EZ%�~���^�?a r���+Y��=�5�xlæz5_o���ы�i@T��v��ŢŲJ1ȸ�ĿQ,��L�$���"�K�[��ۮ�fJ��yv��y�E1g�F-ި
b�P�^ɳ�$��!��#����c�������K�l�Q��29�)
8��O���m�\��!�>���)�����W����3l���I������t�&�r�1�i�l��̘Y����L$�#$�a�\ �o� ��zQ>���l�}�r����Cn�P�s<�K��{��NA�\"N%r:#$_3H�'�J)A��2c1�a�C�^�p���m�Sꂡ�W�/���w��ù)��#�A����Ӫ46�t���s�Z�z`�G�����£bk�q* vg{��� V��Y���+�o��pd�y��1pV�����@V?�4��ܲ�]Y�|DF��\��<��m5FM�֤r���3�9��QL�z���-<�FƒR-��l'�F��Es�vh%hJ�5�}��
��q1��T�E!���g\����p@i�;���d�)۫x��L��1�\�]J&��~�w�0�_��=!M16��r0_]����;Ie|/��2��9ͪZ�x�U���]`TѦ�FϤ�7'�s���a�b�:��2\�X�z�Y,5VM�`/�V��D:Y�;����E�õV;�	޺�O �m�aq�����<QdQ���a�|9Wxa���nv��*�:{6�$�mB�����
�F�[�CP,�U��mIl����ݐ�������삞NA�+�lT���G�����8�v��DD�O��r��tQ��?�����V-j����f��UĽ*��*�pO�\�\�EvO*@��g���"���t�Ĕ�l�y�V�!nC��w������>RޘʟR�@fN��3 S69olz�6Q��E�Ga��"L�������O�P�GĤ-�U�5+q2��|+2�j�NpL(�ǹv�8�l����c��ºlKdb���#zg� j�����Y��.T)r^����D'�✖�v�e�
wƿ��
v��b����&+ Kb��Ѷ�Ӌe�E5����p� f�uS?֌��/Pgm�h�i�H*=9��Rg��e*s��/5���Еt·���5i$�T�a�t�_�Tb��e�o3�n�p�]{��{K/�g�KI��I���������8?uv	������%���jI�B;h��`n�T<��P�"��;#e2�ή"���ֱ~�U����Sc�r7Ŕ�J�ԭT���.���H��.O���ɁO�^��O"�V9�_��f-h�F\�jH��yԿ�A��!b�̧�� wk�a��U���댄|���]n���rx,�2HX�	�K��sH���Tf,6[S�X�ͺ�Ms�m��������`���$��5bB�ݡ����+P,P�͝ �v�o�s*��rS}F����>%�鏥������.��Z�`j窄H�$�LA�L\[�TG*>�\Y��,�-��,^�t���<o4�%@0P^�������6<�V卋��]X�-�ep�aMI_��:id�S�s#����c��o-.k�D����������r�1j���I1E��TRs4?�;Bd�8���	೯����b$7h��û�ְ�6&�[}0U�`�ΘH�b�op���M�gW�^D�~a9_xɔ��Dx�c����(p"�[�g���Jtay�J����B��H�U y�>P�!��#�/���r6�x�F��o���ݜ��2�H":/]�A�T�P'�\D��)Xx S.d�+V=��,���V�P �)��Q�n�m qqi�C�e]L_���3J*	|�x2����/6����$ENG��#h���zP���!�p�u{g��)�P=��6XT�S#�!��(s=�8^��ؒz� e>���Y�?�!��2��JU����٨#�l��ʿ
��Ph]�5����K��p�I��L��G^Bl��n��#��;�Nȥ��2�g�e�L�p��w?�{�:~3����m_�4�5����o���/�~�9�F��L�_����|����fA����.1�eB,sG8�"�Ǻ���۹ǖ2\^�y5���G��i�~�`ʲIR�9�C�9i�"�_�G��T��TkQ�fY�)�wl�s~�rS�}ɂ�������z�� �����zcl�C��,R:��7�vX���0��$��в�����K�5�/[k�y�/͐����*���°nҗ��0�,?B�z�������k��Ms�����%l�[j�4B!ưuQ90Jh�,�2��\n��Oѽc0�O~�ˋ����-��*84_����H*��o���p�8PYfG��Q��C\�{����C�&'�}��:�Y��1���c�bZ�>������}����G����a�Z����=����x)/r�]���@�s6P�9�<5�-:���"�\�vi�&YO��QԼҪ��!�>!�r)i40>`/�*]�Q9���O�L�?�V��㽳��u�ͫ���=���ʫ6 'M���P�rOb���B���9n�p�w�o�ߴS0��$r��}j�R�-��KI���:X��b��b�����:~��&'@Q L���Z�knA��{ʷnE�z\))�����ͯO��wm�)ۿ <E��*�D�xW����I�����G�"�	����#�e<��c�O8F�T�ᩞ�~�Z�*��؎��Z٠�ʐ/�~ڄ���N���f��#L�/
�ֶ��a��9�s��W����_�[������acś� �Yl���P�t�W����6��J�;xjG =�B�H�7�x���-�V�	_QW�>�-6��������e\r����:�C����f����D����g8˧l�1�J�}����k���L��1t������ڑ��}�J_XT�<i�������LXi���o��>Ϭ�h��%]�ۛ�,@�C�E�tfU�b��@c�� �k�6=ڝuM�Sϼ�F��۩r�uغNV����(����狎
�13�S��eto݁-���c�'Hd�I}R�+��'��������VS�A��gL|�`�}n�'i����J���-�F4ሾ1/
�>WEL4\�̬�F`���q��&r-����m�]W���Q,���"��*���G<	�tS���8�Y�y
$GxOnF�_ag��+�P5jF��%�d�]�E��B-$�W���Y�k&�n�*�\���?�<�ϔ�[�)�ۅ��b���"��n"�	zhV��Nm�W��_���s =$nL����j��@ck� ����kF��L�6����E�]�����1Mp�Y��C�m�`��1�#�'6DH�(H=���
��m�,H� ��h`m��
P��p�?�4T�&�u�����Q�9����?��ǫ �'����2�_잒Щ�
C�y}�8�D) �I{�׹
�E6 ����[7�\�!W�V����L���ʩ�>-#����9��/��XB7k��m�����T?�U�z���v����]q8�����:�S�莏���lF�V�]$ʁʇ�&|d�K����Lј�w����ݘ��;w�B�_t��ρ�!Y���-�؊w�<6��m�q�1�K�ál�i?�����a��/O�|b�'�7�2g2(	J#�B�L/$���ĳVC��W��_Aq˧����y+]f�R(3����!������)z��v�`G.GN_����]zՍ\�b�ᚴo(�>��N����d�i�mQ�R5	��}S�������}����^3�p8*����P��TD�-6Bv4ZR�=ն;V��P3ֱR��*S�	��_/�0��,s��a?a	�i��	���c؝��Q�p��2��^��PDh�؝�t�[���J��U7��M��cei](������LI��4�VS�����M��~A�V��=�y`��$��􍸿���J(�G�v�[��w1�S�Y&�i�mVH�;���_��\:5b�M2��؁�����j53����,o������x�mU�'���G�����QY~���_��G�\@V��\�"-P�+H[e��@�+fB?��<�i�ヂ|�4�wN�y|���������cnގ�lV���Qk���0g�P�y��Q�?'���ER��[�n��J�m��z�U�3뾂F����{`����t���h{Avn �-��o5,jb�ȧ �#��Gw���l�Bg���	;��18�rW����F���3��azź�?�-/Ӳݵy������wڢB�g�r6��8$l4d�l�s���v�k�9l�Z��#���Ƭ���EEE�a1��'%"S�P��і�aҴ�r�;9��A�^�E� �a����ޫoH��gѩQ�:�)�x_Q9���<�
14��,N}��>�I��+���YNP��zm�M�[ڑ��<����\�ň��$��"UU�_��x� �EL.�`�y��+������d᧔+oi��c�2%/|(��Ul��O���N�FK�ƐK�4*#�׾!�a����li4N���A�
�)o�>u�&��ٜ�c+��o'�$�g1�k2�+O�\J�Q��ǘ�B$�sO՗r2�ڵ@�X3|�%�uHj��"8���z�i�F&"�9��	n��PN����'%��9дm�LĂ�h�`~ոТ���|N�VUȨ�h;�<X<�*�[�=^��a�BPQ����4U�L�6in��C�&���Fk^��.}@,w4����H��9��Ă�����������@�Md-�c�5`$e  �!���|릺�=%"#U&O�q���R��̖�����B����Qv,m(1�*��L"`$�Nqe�V��;�&2�{"/J@^DOɲ�Ě�'{߃W8�O�߂������Z�^�5u60�zGz�a��D��VX�J����xm9%���0�^3��}�D��q�:f�U0����`��#E`8 w����ݛ�z��mZ���	wYE�P�꼍]#F��x*'��E.�xi�V!�A�=���S�Rʉ.٩
�X�,h0�=-��ϝg�bPs��E0T��U�)��n���MwS��H�0���,8Vꠠ�{7x zz��v��G�Aӄ-Ւ*�YJ�����[��P��[^�ʠ :C�8��;Et 5��{��wK����H0q�G�6,�nX��$3���~L�j�o�f�*(h{�:�z;Z�H����J�z^�gK���8��"'� F����İ����P{!gM��N+��j�u��7�\%�ќ+C�������J�p�F�ݛkf��w���=��A9IH�q���EmQ9�>��-L��2Ҏ��.9p�^���0����箥*g~IeL�
�;;Ⅺ�A��@tlR1�5�&����>H���e[ag����I���b�mDN��Ƽ��f�GR ��C��j���M����
aŵ/k�yY���ɋ4�8<�~�ZI�,2�K~�b�s+f�E��e;|�A4�<�R(P��\�h�:G��k���P߯h��JF��w5l@�~ӽ�eN?�3'Y3��Y�ǅ��b����d�F��I�m��:9|�V.�Z`���J��;�`c��z ���x"ֵ~�)����E����t5w�����7��Uq�с�k�c�H�C���6�T
״�E��2� e�bG����'�U�I�-Ny������*O�q�q��}A�����/6�;�6$@*�0��X�\�4�������?H	c���p�+��n`Q\�xk�m�W��0 ���.�C)<j���᧢� vQ���P�Z:p�b�#S�q�ѥ9��L�V�Vh�-6����-e9a�z��:>��>x���{��K{��}�k���4�P^��[X��Ӆ�g[߇���V�1��3ӉR���� d��$�9/\�Pߏ�=In�S|L?[FN�f��4�N1���j�wK0�&I�&�Ѩ��*��Q�Zv]��]%�',A�l���t�.�d��AX�����S2����9d��KnN-�}������-{�~�a-:��-J��zjr��\Yp�I�,*?���:Z$v�O�9[a,0��ξ#[�Kξ��6)�t$�0����<��,�՛~�
@�o9
�c�H6�ݣ��{mq%�8:�1�T�k�;j�!�O@��[j;��������
Ǧ��v`��k)�R�.?���4���&[_�|�ܯ#!�co"��Q���4��Ѿ1���̕�I6��LQ3�g_�l��A���i��UD��Պ��`D�|k�򓤊�E����#��m�'Ah�3��K�0G�D�%gـh��W%���mvn����|��6���J��"�|���l�4�w�������!��y�Mi���*e��en����E���IݕV���/}�^���V^߻��^�l���Ƹ�ea^�r��nrK�|��r���l�s�.���&����0�w��㶂̤��w�*�����`�ˊ����|�z ��6Ы� QN�����}MΊd�BJfM�~������X�R�\IEzSеa6����jO��~�L�E�錮����6ݺ�0��%TŃ�@��X·�9�·�U٧?�ąd�
�It>��Dڄ�W�'��pRq����gv�ٵ�x���M���JW��c���Ƨ��yh���7n�M�yx��7�Z�x��2�b���5l8i���������~�)F0��x΢���}YGzfT���Q���w�f*�̨���οg~�5��f�\���R�Ĝ�ꏫ(^\���x��[����(�س%6̉R���3���5��U�H��d�y�-G"�?���/�VoIW:��\��_#H��D0=��\bS��3q����qY��}|_!�rM�Z�@�Fʒ-�-כ���R%RNaqa�7f�Y���^"�e��C��$��$F񥚣�U(ɏ��P�m~{	;~���ꭍZ����Es|H�FG���``9������{,���2�%��"�!ǾQ���'�U~<���^��%mݳ'8��&EzТ����d��Y���S6g��w��'|��41�N�K�ν%���a���ՠ΄����-�p�q����p�#nX𹉁�n��v�C�蜺�k���Z�E1�5i�]�\'�B|Q/�y��ަ�yL�ߧ��P�6�r���2���Bk�9H�#�� ��4������ �JJ_����B�_�1MB���jj�����l��,B(׉S/�]�;������$9^i_�_&��p\���Z�����^��b�� ���7v���@���r4�3�/2�~��33�&��}��}[?�4�e}𗭋���Og�r��h��P��ԽA.џ�� �7#t<q�6m8G��Ι�B}ղ_-f8����^�"�� �g�B3!k�;�$�n�W�ŷ�
�]�d�`|���	�����`��F��	a0���k)���e���q���P�sd�������*������0܅'\�LZ�"��z��J����J���Լ
x�{Ù;s�Jp��IpOD>����3�]�����p��%ceh��6���K��=�c��+��6���$�'#uF����@�r�H��R7?K����2sW��Xw��C;��x�����=�(FC� :��&��/�*k�N�#)2��v�����;*P�6-�*Ε�-�>��Uom��
9��6��J�o:Ĝ�^(�W�*rMR�}�l�-r�~����$J�Dt�'�~��2lsf�
(KƇ˹�?LvD��t�Ll�*Bu����ۨ�ŀf�'�o~[�'�sa�N\�#�m5A�T�Xw�M�;�F���j#�����*�����X&t���L���������K��J�c�?N5��<�א���D�d9��i5��	/�E���i��l��l�`'穞̿�P�'�~Δ����6׌�*�������Fv�\����E2�U$M{hZ���6C���:2�厚+C�ք�2�M3yIJQ�r,"�0���+7��6��D������"�g��"+��8��\:�ނɛ�@�{;v^���|��aSP�%�e���g��}W���U����_���uI��c"Z�&����j������ΦHBw%�/�X3���j<��4X1W�:�]���p>�XpMF*G}bt�x���}�T���S���%����)x8�H�	��x*;Sb]2�lX�,G1���6ZCz���9�U��?�x�1�=���������P�τ�Tt��o�~&���ʸd+(�qG�&P%�8�s�e�406��I� ��fIVf�L0%�� �9^����XhFY��UV�p|��:U�"^p^�XK���.�޷xM�ľY��6�q��Ъft�'my݀j+_��"H��A?P�Xf�``�^z���`�9U�d`��i�&�8��]9	s����	�����?Ze!���]2��6p��#L����}�J<;P��QY�jZ1'{�)eƊ�˰�*��	���Cb���a�0U�<�0���E���	��7(+���ƩtH��hܦ+»J\���8�s܏L��s�mY����g�~���/���<ͽ�F4'��%��p	���Gs��@b���E����9��E��E/��<�m4���Ʈ*�E2^½'{��C[NA��pnE����J�m8�;썡�H`�A�]�;A������/LΏܪ������\����c/50tZ 1 �*P��kGl,z|��)6�{^_{׽�Ax�j���X�s�����2g�@%��}	g!��?N+XɨV�Ȓɰ�Q�Gw�*��Uۻ�:���f�Oe�^��.ԫ�ph�`/6�)�S2S��11#h#���$	��H�Xl��s��r
���.U����İ���z,���H�":�Lp������[:�J��o���9���Gz�W�UC��E#�l������r�t�Ŏ,�y�T��J)�//&x�4E�� �w�h��)R����b6�},0ذ�\�޶�՞�3�bA��E�&�!�V�g����4��j�^_J�?�U50{��k"+`��~�O�t�����I�H�R)��Ҫ,�І���%Q���_�x��%�1�=��=:�Ȧ�o|jx:�T	[�����O����yU��6�L��%f���%T�*�0?8J�VZK�������#��nq��D���^ꄝ8��{�
��;=���e8S3TfT���h���)è�_�L*��vj"�!֧��uW�(���PjbٱT?=����ש�98�4��^������{_*_�,?ʒ�(���?�+�`$L�'�{�}%���t���`�>��1Ҋ���gZJe>��g2���?>����?�����(ALfN�l�N���&p;h��`[�ȇ`j����'�d�E;��=�����x,Ӧ�1b��魙�T�G����ew��k����0V��pLQ!" j��fOc�����OȺuq���'���ze=g�t��7�t��-��шF:�Q_@�|�(%�D!��X4�雞�nφ]�����1w:ŤD��O��?��E�Ї㽼���|V?�N��Ő�T�
ߙ�	��>���`q���[	7`�H`!p�(� ��I�}�T����|b6MN�ɰ��d�~ʦ��U9���QgD�i**M��gp����&b�ji@ ��X�Mlv�l�k���)�c�U�ܳ���Ͷ�����l��v���$�jH���=���f�L�h�9'�qm����-��{�P��߉�T\ ߞ��Q��~�`���.�C�q�O|�3s
���HM$��5� %��`��w0S������@��L�Z��MH��P3����d�<��HT;�8f}��=��)s
<��=�8Ak,~h�TԅH�r�͟�G�|�]"wc����th��ʵ��r׿�.����Z�_ܠ��@Cgm�Г���};`D6��x+%\��~hC�y����̌��;>H3c�d;�4vT<�q޿Xi��w¡5�} ϖqU���JʭU���2�S`$
��d��d�-�hn�<Mf*��qT@ރA�$jZ�[__1a���N�bj7��9`ˤ���VM�6�B@�6YQ@���r�)�*�TWL�Ƶ��I�}̎I�����F�O*^����1}�����+k7���	a]/Q�go�qL��kI�X�AB�.6	��_�5^sӫ#�4��L�7�&�j�����^e�A���,�=2~D�=?�cg
m)��.B�:{9�m�ie� xd'N���J���Z�%%5Vd��s�G�����;�R��������%�,1�F>����Xu��cv3G�m�	�x�����4��mߡ��x7��r}�܈S6�5��ZF���-�i��ø�#�6D�Z2�����������`�O߮�2���b�\;Lm837�i'?!N��x��	�e�0+NA��� ��\�+q��,m�!u���уi���M�Kb��$T�#I8����ڵ\��{4u�B����t���	��Q��.}��oe~��ӓJ,�[\e���-�'.H
�[��B�ɰ��v�,HpӞ�K�%/2B��Z�X�2�籖�D�G�Rq��ߜ�����Y`t.�mn�I/�qn�Ãq����d�N53�����E�gs<�{�~�6+A�fK��EV`��#)G$~���$\��=���B���,�x
D���~��Mʂ`�܋�����*d_��[S={'����H�`,�p_�&M~�8D<�1�E��2��Eznh6�L�.���#�����ޓhP��L��@ި�� �4Q��K{��G�ל)M�x��BW��I{:�p3Fk_+�Μ ��CZ.A�ʚ3�u`���|;�s#�C#�{�-����N�N�y��f�D��.^�9��۳;-�����T��P�(��t�n�k"�Wε����wo��v��}��ll�9@pvy��WW�B��.�gi0m�P��6�*�Ԧ��M���=���ȷ�[-��.�{�L�8Ѽj.t��n:+�a���Ƶ.ȟ�d۟[���£M@�%+�rr8d%���2��]�����'�2׈��'���, p8��A��u���M4Bf��q)Xq_���;����gbGhH��L�C�̰������`��PMf�]u���\."��?���f7ƴ��^*s�}K���>�m�* {�6��l'|��v-���DK�Ht�g��4ZR���|� ��@*���F|K�X��%���1O"��
�NҊM�ؤ{����{_5��f�Lh��rg+�?�#fB�J޴U�%5�.�g�v$������X9�_v��T�屧��u�F����t�@U�*6x7��W�Гw	5���(=e���w:uI�mޖ���U<I���ʂ��;_��"� ��|C�����B����5�b�{�N��;���`P-f\�[+��Z��%�� b+Q�<b�%�u�[OKE�9��q��;j
��;fR�s��@��'� &�(1!R�E�,|�7q�R�mu��(��� � 3�-"�`Yp�8k�k"����������|N-���`h[=Ø�A��"�QPs����|Z�?��^���ʑ�7������H����"9aO�l�۠�5,��@��Bp*m�k�1����-�]*��������_dRֿq�я
�Հv(g��ȉßZ�~��[��V%h`ŧ~�W�L�X5�;K��z���LbXn�*]UŌ_7���f�Ԓ{�h��Sn��P)���lj��N�@��I~�3�R�;�L�Q��Ӽ���+קS�'�)Y���X ����~OEHɍ�҇�����`���s������'�E����ry�����TʔJܞ	k+�}�=��B��k.�ɕ7�{�$�ҽ��x��e�>�>qV+^{Ⱦ�ę�5df�&���㫾��z2:id���-���OUd�LZ霝���*�g�]x�?`Hj�5Fi�����p3n�}�S=�?F�����؆Mͅ���� og5�Ïw�����&,ȩ�&x�{H�aQ~��6�bE=3�,��W�ؿ��I�xG=z���g�+'�b�r⽢��5�/o��\y����H�R]G�)~X{qeto�{��[#�0�������p-�v���L���
��]��Q3����W��(ḰRf.�812J��G5�ʀв4|^&�۴?�N&���@`.��b�<�n"���ڒ�k�5��oP��K ��?���!������4�!��/�_��P�2�m��
��z�����1����A�c�M_��u敏�S԰��~"�}�����	 ��ÄBi�
��7yIK/f�"�O�aG���Y6�X�2��:�ڄT ���[��9���Q��@�&�����z��3~/�]�{��A��iC"��d�  ����\�D��[�f� V
�ď�{���R0u	U�_�x��̥:�9�!��E�J2n]��	��O�`�P(Y��g����H�����6���B�b�m�j��<���-��1\��c-�2��C�Lԁ!��|�Jt�C�=�9T`l.0�<�S���Z�˹�R��;��v���N���Pf~Z�C�Y��8���NG�J���?+�>3v/�o�GM��2�~_��?�֗���7�o̊��y
fo%sC�<�J�����>{�d&�H�#˄�ȱA�q%EO��ɟp?w������@e��'C	0F���t �P�g�t�+p�t��9@^�B���ʜA��x�Ű��QݾA�M�g��b=4��a��}!i��jH%nb��:kd唃�il �@���W��(&�ȅ�5�"���
��r�\��ߺÒ�	>������3�B�e]q�1ѝ�����iF����ۨ��nao|�	��c�,1��\��C�������N�q��T�ƥ]��?i�h��[U�D��7j^�B���n>j=s��vY9���p4��[�"�vO�UH�9��4�A��'O�=�8GA��s@]#I�x�
>G0��{6���M��[�����6�[��[oU��)S���S�"� �+j(�Z�?٥�:��
]V{��@S��,�����_6�ۙ�j��o�]
;�ה��EV� ���>oy�ut�iD��� ����$�{0�+9�8l��8��د����`q�Z͗ͽH����eWS-�s���r����fL�D��{�R����7l~ ;DP�ǽ<\�T�jy�k3�l��%���z��1w4��i�pS_ɭ1�$ ;/��;�F��y8S�V`H�����j LA��4G��~9��G�V(��3z���*s�1<'���f_��r�	�ch��<�e��0�� �R�BY��6b�7��X�(��W?G�B�b��A5x�|�̊�!����(�W�'��bf��Vu�h� %��G��*��&,0���P��)I�<��xég:�d�Ot�p!�Q����ֺ�t��$*��SL�p���Ĝ��6����Z��5"�|�R{�Rt��B��/E^�{��X4�c	F�5�*8[8�ƞ�e�`��A����j���2E1�F����Z0�P��4"�x�A���̾-@L3a½��5fb��}��ȕ��/�M>�kG���;ˌ�-�-�}�G�t�j��h�ϭ�m9��RU�������|az�0E�z�(~��p��I�q�����T��G�v},�����[�J�{�1�<o��@��D��a0������R9�U�Iƽ�np�l�aY��Z��{&��"U��q���H��/�u� uŏ�WE'���Շ��9�*yE�k0<��>R��D̚q��p�)D"H�@W��
ƍ��$��Ú3q� ���Ce���T����S'?ޥ~��m���(�gs�|׿������E+��BT�}m��&�s�����*�����j��Fu�������9�%��N~���Cuc�`cje��R_̻f�v:�a��6�b�� �2a�/r?`}fKV-#z�)��YJa�v5��#c��@+����C\ȻV��!A��Ul���J�kD�;񿴕в7��2���������5�����?�,�m'��ZK��-o�=�����u��p���3KH���[�����:�㪎��"�TiA,�����S(�h������Ѐysb��ZB���r���s@s������r	Z5E���=BO�J�፿.��_�jQz��N�C���)XI�un�ެ@2y���1>��@o��C��CsbŇ<�]�FӬ��2\So> }ԤCVv�� ����+Z��y�Pd�������&�r��#F�<#��)�-%~5/$|v�"4��Ƥ"{^67c�?�H� ����0��_��AU���L>>W;S���A�x~^��f1I�񅰮IA��	P���6��y��Jٶ�$z�٨qY�:�N���t��/UVyn6G�}9���s�"�|Ӑ�� ׍3��za?��z�T���E�M�?mAr�!+��h���2Y5)gJ�ϖ��R^*##�.66���M�x�j;�m�U��NG]d�	8�$p���!�l����o���M���>�ݱ9l����ّ	��e-���;�i	��Me��k[�����y�I���@��)�_�n)Y{���C��Se�D:SP
jgY��
���G��1h�+�/���J
�[���%�ea+8�rA+͍� �B��u[Y�^�@����-�+�,�u׌�y�����:�|��Ec��97��W7��0(J�sgr��q�X��!���ᇻ����'N��'�:M�@Kڢ�C��sH�]���a��u�jN���0�F}�o��11��(�>b,S�J�~i�.C�6^B���7:��̦���n�;;�i��C%�,$Éd��/:�4r�HԔ�����,������T���G��ISKۨ~Hb���U���� �Q�h�4���4��GSw��3�h���j�	$��0�ܥ�݇�V���r��z��A���{���dP�\��ɝ@Ff��&Sx�SN�@y���C�c�����T��Ǳ���k�k��j6S��c"�`ۣ��VH��o��MI_�K�wi�"ouRґ��a�U����3��cn_�Ղm�k^"��<�00
�y�\a<�]�lA��t�n��b�o�Lٮ�I��MR��.2\��wi��"̫"n#�I��IZ�{�]���Y�b������h��p?��n���8j��3����W��37��)�]8��t�dh	K�h��G�[��J�}ɀ�/얶O���'�u4��7@��Ԛ�Mר>,�NQ
�����Q3�+�*�ڌ�G�	�׬!�u���4�H!t��>=�Vh::�{\��h���T���@?�cQp�8I�$p�����v����K�zr�\:�f��ρ�ZK��������`�G����j�f �f��M�i�gf|�wtSp���~�Y\,?o��r$�p�M���˿Я/�:�L"������fY��{chA�M�H�o�'����m<4Hi6�k�z��֕�x�:�j����;��Jv��pǙ1�q��8Z�q`e���$_<�L���,�Д�P�UY�Ag�=?K���NtÄ4�	�{��.ݶښ�B���9[Q��ړ��/�#h���k�܊��u�} ~)��z�87���=U����yʒ����Q�� e�r2=��U��쎔<� @x7�c4��-}���U�DT�JA��߽�y�E�����DfC��j�P�����O^U����IH	���L�wr���.ȫ����M�b!y��3���K5N��Y�y(��:��#�VN�R7��b ��]�� �Y�Ԙ��N��B�242u��p�K@��u1����u��
I,�r�4��K�o�$��j'�;�?�L�^���+!+=��7���B܇:C:l?#5�:xI]#X�_�^a�g��Sy���w �v)vk�yZ�4`߼�L�>i'���&�'��u%vZ�b����-S�(k� �"G\��E�e���]�1��M��^c�]��Y#ϗ��s9/n*�,7Q�'�L(
��Vg��ѳ�,��>�R�����ZlbrH�Ϯ%����H���	��Z��2u��*������Դ�G�«LK�K���79�DD�9��3݃�0*��k��l�l�h�86�u!k�g�u���i�EK�Y��Y�P��5t]%��i�Z�?U�N�ռ!.:y�sh���H�'�B�,��܉5(�ٚ	:�!��yG��j_�u	ٸ��iM�g.��m�����b7N��N�S6�hgρ�p���9gW��0�]&��&�t7-:��֙$[�㦒ڢٳt��^�ǨW��Y1wf�C��\�SWb���5��x`Q	B(��kfX��͍���Φln��Q��v�NT;x"�a��6�5ejS�@#�FUUm�%7��e*B��c�2��~mW��#�؁3�)A0%�E�R/�'��bJ?^R��P�c�6A7�s�\�<4z|�uKW��nG��c��i�m�i�i<ƭ����L�x_�"���b	G|WO{Ʊ��ؑE��BI�\�ҷ,�-ٮ�I�����!g�%�)�"j�[/�ŲEƖ��u�$�w�u[���f5�1�B��9�+��i���b�m�qo�i��;�O�k��ZC ���N}�?׋�27����OHR	eM�U�
U^r^K#��E�0�� D׷:��s�ZQ�mC[�l>��U�8ƾ*����)o����F�\�(s�"C�޽� �2�E0�l6�,���W���c�������X�9��ϩGcJI�e�n02\e�Y+8/�vkwS-�3=s���)v����b��W1)���5S5L��ao�u��x�3�W`��D�Ƀ�!�2<�>�&��x_���Dim�rN�	JK��8j�
�n,�G|iF �KN��z�ը��눹��/��w����-9���͛��̩]x���KS���8ђDT!�|��ro��)M�c�,��~n&�!�c�>��ު��	߼��T�lKT�!���c59\��N�nN/_};����yrK]I��wi>��^ǻ"A�4]�[k���G� Jl'Y�L��zA��ŧd���
;��t��D'��H2�y��V��~޺C�z��PH`la������ϐ��ܓ���Yy�zd�d4�	R	;bgة���� \<�?.�!p	5'�\�H��^���8&��� c�v��
�Ǉät���ba3*1'!�1ث�4���h���*{��+Ob+�s�h�t�'@t�/�H��W�bۧ!OC�*�L�ˑ��_fxYF�"({��/5�����	3�v��jlg�m�s��ZaX:X�h?^�=��n����ؤ���7|�&�,@p���J!F��T�wc�P�N��t{*	�#�;�mvf��N4�����Ek�䦶��07 ��{6��'��E�;�W�l�7@d1j�ٚ�a�`����°��I���)��Ms�>G��߰�+�YR��I%�Q-fԝo���K/��b63���I� $���:`����Q�� Y �U�<�,��_���N��4G��Ob���?�����>�����n���@�)F淳�x��t��1:�]�Ђe �-�Q���Kz�����,�� l�r@���*xq�Xبn�2�m^�k��--��/|Op�/<��O�P�f�anu�ͰWr���ˢ�,iz����W�����	%����rU-���e�񱡔�-a����@�����w���p�#=��vǺ�DO��R�1ԃb����qK_#j��|X��å�l�u>%��!S��/:Iq ���S&-l�y8e8,Ͻ|���F`L?�M��Z�ߥFVB�s�c�љ�!�%�$����T��X��"��I�m�92�`%���K�(�|!f�`E��2��z���X50ge<:Uh�tOY�Ǩ#��\r]G[�?XMA�WVzb�M���Z��΍ݮ�F|�L��Ӏ�ݎ�M��{�r�+�i�s�����Yt°�wȲST����pI�6�X{d��H�A�<4_b�OЍg�����cf�k��)�)9�2O��=��\�y�c�qof�^8��N؀��E��Vin#�9���}@l��C�i�~�3K�n�Q�	�t�Y�ؘt�[�G�~�%�Ґ�V�f��
!�Ԕq����zk#�z*BY�W�lu����/���O����k�UM[�hy�C����o*��6���O��} 0O� oا͡��jEC���k˲)x%������ԑJ`����2��R�ȇ�Iģs���t6w��g2��_���S=�j�c/�v͐��H�����r\���䴭1�ߟ�ޠ�pg!��I\�2���ּ�ݯn�^k�ex��VC��Bd��mɍ�퇮v�-zʓr���רC-�� ���T��{��:ǚ��y���r��8R+\�qJ�=����4�a�h�� e]H�c��X�N��M^s��U���K��^���w�
�7Ù���xg5XBq�X��"!�519���X2�7�����?]��j�ǫ��Ȧ[��-U�'d�_�N!���K� ���Z���ʗ��~@&R�D���9�%��l��G�������ɻ\v_zT��,�*��=��^���Qå��Z���W�%Ay��E5v��%�2��}!uHlY����E�mn2�Y�Nϛ@�"8�x�^�:����'��N���5�q�#ި�T"bhr�v�+��a�����!��m�D#�y�s���x�0$ߑeq`�^���]ߋ&�%6�U�=�2D���8p���QKEɠ�fFƀ���|k͠wr�X�����ȹB�B�Ժ���2W\y�_M��M*�S�$�t�(��*�E�OC,N�4��6�B֏jڏ�P��}�P��_%��C�%LX+�G���
��Z��Wb�)�7��t�R=J�ږW�f'(>������q�]�z ��_�1� ��8�,ٝ1�8�ː���i!'hh�G!�|�bT>g80�a}@R�dk�?hQhGzW�6>�m�40��*��0����e���R����	�4�_���*�?��՗���{���3#�b��wM�1>��mDf�4g�I�{=��^�~2��r%idp��Z�*y;h}���
�n��,��V�b���@<TX���N}\�)�����9�k���А$d��y,��"��m�E��+9D���v�$� 	G��N4u;PZ�z\�@�y�б^�&�X��|o��|��6C�ᧈ�c�:*3�\�\�~��B.�+jCi��|p1uv��k 	��X�t�/R*��>��5�Ҏ�W�n�5�0䧽��{W+�p�A��ɻ�ude�R�p��PB�YK��j�V����v��{6:7�-&to����w
�Geq:�!�W}��z��g2��u��^n���o�.�Uirw���T,�Ū�����etV#���
/��u��R�2'�����h� �7���G�V�%�  vTg��.(bj�=dRY)ؑ��n{+��U��z2�<�f�|����ڇ���jFN��H����#aЦ�T�đlp§�afb[�-^2��a~
5�L�PM{�6ǂs��?����������p�{�FA�\aʐ;990&����1�=�u��O�؎�Fέ\��c��6�����A�Y��7u���yl"��N�u��9��P��O�8{�DZ�+#�4P뻜���Z6����];�D�YO�d+��*��í����M�� ��b ���ݟ^�|𢩍v/\C�'��.>5%=3��kW���%=���:,��6��a���$���r�_����/}�_�pq�#�uR�=Fu�����2H�8+4���	��^rk?M��1���ם�L٥7Buo���$���a�Tn��:!�N��vZv�����q�z�V�<�("�8��Op�x��b���O���*��Q^�#��As��`�\@�.��SCmH��z��+r�/�@��☀e4�	�䏐1��I+�����]���SGe4c **�bc
��d�����{�+ձx_�����=�ѣ�~���>m
oQb��٨a>\xA��7^m�����#nn�z�����n�����)s��K��P͐���v}�^ں�b0c��℥�[�h.��-������0�|�I����u����8,ւ�oEJ��z�I�/�D�D=c������/��lm5�h6�om]ް*��,�X��E��@�0Vʻ�F���00����nFO�(�nz6��V����{_��5j�F���Î�@�_ ����>�>K�*�Mr'�{��p��t� ���˳�B|�:�a�2�P�O�ξ.��_��疸�� X���	(���C�;N���i����ݡ�a+��:�|�#�\@�c\��=�?�|���s�.����KK�¸d�2��k/�n+޳�T+ޫq���4�x]R
������|���Gt�ȝߑ���J�L �<��ҚQ��Ý�;����)�|֗,/P�]/j�:�����,"�V9�巐}���+x�����Sv!@��u�QIA�(t3+R����˞����������8S.-2�#�X��7�7Qd(�P�6��!�=ۮg!r%�-������ɠr�?�tݙ���NN��áA�I{u ���z�����۹�"<sZ%������_K��cS���-����a�[���0R��#z��J�������u��ɣ�;�~2���m��|�wmA��`�]�lP�6�� i5��	�Ce���c{!���[�K�y� �ڌ�ē�t���1�J�GCՄ#�pR���z~xA�"T�*P�J�I��-�>ª� x}�	�E�1=.p퉼SD�Ajt�[q?�n�HC�%�w`�׃=����߯8��
�����oh{�b�n��QQY��a�`�Z6�i�����W��=G��{�|Y{ �3�<��"�9W<S�����0�tdą�p�:W�ep�O�Ќ?A���:�d^?0����~�^� t�OC'���\�� l��S �+f�ӣ#S�B�n���������h�+X�M��iY�̍��U+��]8e�f�O��3���2K�Ÿ��sHjU&z�U�Eє�0
lg��敊+?�����n����6eN���������HJ
^��s:�3W�2�����3��{��è�ņ���I�+�N��W��}f�#� �Z�B��J���~�� Νh��?�d��_�8h�T����#��r�t��~ >������N}1�+����kԈ�������n��2R��6v������ͽs��7Ó�B�5r��oS����̟�9���!�s�)9ክ)&�1��-�ju�<#�z��`���%�92���{�Q�i+2�$��! qye]N��v�5_D��OQv-�t�AU�`�N�2Pz�5`�@��ub�s��w2��mX�[4Gh��B1	xB��vs̢e&����ɑa�jJ{���&��-?2,q��q(��|�,q5�/��h�3Ԏ�E�R/�k��f,>tqCJKO�f� �����(q�����bj.��9���k����?���+a�it�)B�9]���)����x�wp��!-��bq�+%����uƟ�Z�Ŀ4f�s�т`%�����'�ES�� ��p��5�����`t�d�녯M!��y�Ԝ�����pk�Fg��9C`�yi��]���|s������FUZ�v��[��b��m�O���]����m���8�|
��"�^F_��x�6��2'�[����/��N��.4�m)Fzn5�:�#�0z.�Oe�1��{$�<t��"J�y��?TԌ�\=��������5 ��~�լ�l�K v������6c\�ŀ����/R��WErT�]�E��.Դԃ8�u"��+��?Rz��6��k
v�ڂ�B����1R\~Q"�ކ�c�B]�G��1����ow���m|��kvxٷRZ��酯=d���)��1Y���EG�<C�0l�t���u�K�A�.ZB��'EB�˨�ov�K��G�8��A��{��!^�.����}ƻC�Q�E4�x^pǳ�*�>v� �`�	�!���R��dr��#r)�S�f༱��ޚH��ꊈKi7B��-�f�ʹ�8G\R�>�+ڐ�s5�Ѧx��|.Xj.L�u"`&�]"���-��cfT��=.�A9@ڤ�B��N�?:�Y^���|03f=8����08	\b��M��e���u�b|��z���,s~��k!`�2:8���Kzh ���*���K���ъkʁ��+�=�-����4�h�u�|�st�,x�:��b>5.�VP�������q��f��uy1���h���0*�h��$7�@��2��:t.G�X�߭���|�X)�x�ʸ�k� D3����Y-$$�������{����16z����w�3�f��g�j福d0�a��x�7_5�Z:��Y[sQ�3�m���މ�4>������H.����zzR�a
��j�GO��`×�Z�����.�{�[d|�8�3�r���A�%��s�H�~�Z�1�q���J��ɚ�/켉�'�U����w�;�QA����f]��>@r�	F����]�蟿�I9�O�C˲�i�����Ky���u (]}��^N}��FD��3�*�C(A�P޳�P��D ���"�|��.pk�<�l��Q���(W��E袌G=�i�L]�^����,O(�M��P�?���7@��N�#��^@޴��z�[3�y�"�&:��в������y���C�_��BX������
�"yw���%��`��Gy���rO�66�p��c�֡��P� <,�%M�n�3����f��z%}D~��u=��բ�a�A}��tSҳ�~78��h��=]Y�as�a2UK��;�:/l�H���Aޯ7���3l�j�SןQ���b�y8��@�X��y(tTiϵ9�]��t�Ƹ�_�jW���<H����Spb �^�kS&3?9.�a1��}��Q"ԡ�0�G�h�=y'2�ڪ�
����spv��x�w���	���S~X잦�2)�?�$l�Y$�B�T�вwa���D�����w�W��=�1|<�a��K��=$��=T�����q�d/����+��k��[>p���S�%�G�jښ��x����;�O����s��uڅ���0}f_�d��Q>���4�rR�#}���;��������=�0"Y�B3��.)�#}9�d]) ?'b�m�!��➡�x}F�zQ�]�/Uv�ǵ�y",�f��͸M��>�M��4�SI�Sw�<��w:\8�b���S)'��9.$/�xF�He�>Y[&[u�)f��H4�,�����J�s/��"���6���?o�ά?~ؤ�	;7~��Ӱ��e�W�S`.�boQ�A��$K�(�7d�S,�ɵR�"�F�����yk]9ok@}G��2�!���in�$f�x
���Y�����YHGo.�#�<���I܃����R�7)ka�������g���(";�̈́Rj�o�����z>tG)!8>�ӓA�ӥV�I!���D������ �ە�����I"ĵ��0!���,of��\ �:�6�Y���W�:���b��X� fb�ӭ ��5H�Xb!����$�N�8�ɇ2ޥ��cBc��5��mE�o5��%�Ull���!W}W�~�MV���F@����IyL4鎏&I�*��X�]�����xcS��G��.
K���� Ɖ_����X�o@�����3%�;�Ġ����v����w�&���v3Gn���H���.(RU
L�#̩��Yba��3H0kRꡃ�l� ����TS�q.��O�|�{N�"���oi�:*�G �B?��[Q��K����';�ۚ4#Ը�����[ZW���?����̄6�Ww�3/���B7�y6�����c��Lx}w�8�r.�)�N�q����Yؖ<�j}�G���=��\1��q���/
�J;��>�11�0W��8�l!��%.��<gs"���sb����P>cY�s(��થ���]�7��vՙ(���<���e�s�S����$��APK�������0��BC�d�>�N��2��z�
W�'�,8$�����zo����
�+�h����kۊ�ΐ	_6�i{W[a	�'b+C%+�$�>��p7/���_�r�6t�,�+�$�����Ez��!���%��i�F}��xʍ�z�J<��)w=L�^<[a#<PX�PT��"pgZ��H��<3�5����. �lD���w�����ʂ������C��A*�=����Ԡv����r<���@ ��9����s�U]T��Jҫ�: {�*,��a^*�SQ��h�괇|����OB����I�>���̝�AӒhr�YEc��;  �aD<u_f��Sǃ��c��x&_>�k-�\��K�I��ǀ��.��h.	����r�Hd!@P͈�#��ioڦ���,�����%~U���D�*�B*d��B�j�ܰ��}�	
3���O�[�|;6�YIv�9��|p��?^�T����;��@�~s/�_D�7�S0:3���O5v�Q)��v�oIS2yDi;u/v�W�O�!jD՚t�S��Р�M���W6Mi�i��y����U�%�4�s�NB/4���gQMd��i��k�6���6	>�.נ��HS�����Q̨�Yv�BkE�Y�&���.�:�2d��NI����w&B��[���&l�*��" �Ҍ�O���k{.�6r���D�z
��1DbZ�o�?�@�R��6=aQ��uL���<Bp�'�����B�X�X��zjH���? �r�b�M&��h�/�u�<c;@?��mL����>�:���]Wy-@��ԘC3y����98����H��S�['�ɣ ��+�5�1�!���!qz�䩸as�.���>ʴ5&z�"��\��0���j��:��gL~�#C��i�N����~F�+�ե&|�`�@���q���ͻ�Ɓb�s�I����I�� *��z�����0��4��#���,b��%�ZՑ�xĿ�����j"�Q@�#5����$�-�da�.)1�[�Χw��w�L� a���I6Ա��o�I娗xhLf�ĳ�Ӵ�8闢�Y�!١뾻jT�8P���1o-�v.�/���*�i2����N0�{˚��rG���S�G7�c����1�M�d�mNUJ�j�5,mF�H��-�V�GH�׈����|g���$����C/zż\*W��"�t*1���k��l�?�A��U�il1;D�?-h1�H��6JꋲO��rDn�R�=^N�؊iɶ�y[쭔"��$l�)̈́6ݾ�X�s�� m?;؃L)4\�&�eԙ���~ Cwn�n#�S��� �^��ͮ�?$\1�[��q���J*���+}(�[Y����e� ������g���,פ2Y+ъ4�mi���0$>��Ig]<��l�&���0��� d���X�B���m��v ���;k���Њ]��0�cT��yhj�O�]��Y����楼��%����6���-no%a���l!4�D�����N�T�U���/]m$����|]��xʮ��n��ɇj��ܹ��N;�q��<Z� v��vf�����f��1CJ�U��|yx|K��Hk���,�'M�Ive��,��� ��ph�dhd��	
�U ����b�6:3RC�k�+.��-�h�uu�����$���󷩸x4� �X���Q�D'H�P�L��iFu���#0Ʒ�!��)�2Y�L�-�}'��v�?��ϟ���954�,{��4,����)��8*��J���L[j�Ԅ=�����q��X\89w2v���2�"��2=t�h*���9K�PF�T�������T�n\��!0MUG���"�����y�T�&�q����8��{{����!|d�fb�^K�c!��,[��s�DB��Y1�I���F��\���E� �|�^ZH���n��g��]�:���R�Jds�}��`�"(vmO}�,�?J����c4*�� �ʣ�|-6e\^�Fη��"UV�~�D�2�zIMu�u���WG�H���O���b��@U?��+����2T�2yT)��J�'h�j+�r�ذ�o�wA�$�ǅgD͝*��G�`�d�h�po�k/y�;�:�؂y�I��a�@�O�F�
4�OS�5�V�a����*j�������͛�Q4�����c�:�C�d��;E��V��6�����Ƭ��{�IOؠ��V.�u������֋JMb
� �˪�~�E/q�,��4� !�E�Tg{�HE1�9��U����߬H�u�Q[u�[���A�6��-3F���,�?�ޞ*�!���>�e@��!n��	�RӘ+L������K ��L�a�螏 ��'{����c��ᰲ�4{�b���}R�8��-���kcܼ�9�Z�p�s�����""��@AM�v�ߝ�oFI���@�lS��������heh����K�˲�]�K��di�]`�r$�#�i��[�e撋����kF󆓴I���m��~ܒ)�,�������}J3�FQ��G���A?�h�|7U�9��/|\�.�ހ^zUE1%�h����Q�JI�7l�5f=�׽��s��\�����/u������K�p�̆:�0ٻ���2�˛��^D0RK����ŭP��XVct�a��r�[�4����!C�<_�v68��N�r7��>"�o<���t����%�Tm�G���Z��X���eI�Ԗ�ʑ&k��4�� LIF�"9���~���1��X��ϸ�*ڊx��[ȉ��tf�LA	��1�J���'���V�ή7�UPG�12��O�b���U��f��F `���ro2��W��U--��84%�Y��?�tԋut �"ur� ��l1�*�Dz&s4�����xf�״\ݟ���	P����� z-,NEEۆ�Ys���c�՚���e�״az�]l��� �cE��H�nQS(zǗAÝ��z�_��*�5�Q�����9sֽ׏}q�O� !�y��$ɒ����|v��̿u&So
Hd:�IJ�Q��*�%g!ؤ����� �QiB�D$�.u���)?�;Q�ѝWjS��b�y�XPg6��8=a�\l���Q�2+�e�I�Vlm�	�d�r'��:{��N��.��HZ����x�֚�XJ���������W��P�a�2��H+C�IV9�c1�D+$��{�X�>��+ۮo=��E�ZGt4��0���?g��#I�+��}Hr�y��j���7�4��%�����Q_�����I�CRu1`�fMQ�s m��g>^7����CBp�́`�$(Ey>*6Ю�<ŝ]5t�y��?�A��ֱD�`F���ts������!��<m���X��v�����E�w�k����@7�ϔ�ar�1���QD3��m�o�u�����AfL�l��s�?�3�S��ʰ�3Q����ڜ������zla�3()aG��_���XLj`�X����6v,X�ޒ�˴V�z("яI��xN�ܺn��VU������)ЁOP���
����)���M���L�S��!O�V��'2�8��aJM`���Z8z�O8�H�Ȓ�>v����l��[¡1��w̺��L�U����� f�Gc�f��#��\ǡ`ڍ���,%0���<_�O��	�Cly�!�n1̚����0g�T/���d���&��=�,������ۍ�ئ���N���������af��5d@10� �����ttA�ti�]"r��}��^"��L�e�䄦Z �m,1�SUG9�"����md"��)�H@u�FV�e�b�7����(�:��i��P��9���i���T:������V6�ʔ0M��A�&�e!���1=���H1ps���(�8�S���آ����1Mo)ä��%D.E|��ާص��J��m6#���:������'29�֖�S�:I|EO��~��H���A=��-Dtsy�ezr��fA�l�o�^�YA��B(_�fA�꘾[���&1����;�H�$��t@#t��g7<�4PaT>r��3�+I�f�ퟓ7�����\o�4!�_c�Ěy�h�Qy���Z�v���
�˥�OP�H}�u���f��iAH��?*7"��_�����A�u,��u+=&(q5-_憯Fz˹�	�Qs�$4��C)�=I�Y�ʎ$�����m�ZN�e\'�…��:a�����iE3�h�k�ah������,�7m���Qp߅5�G��H���1##��Ѵ�f�O�,�/Y�O#l�4^�P��\��ەj�T�S�Wa���BH��Ŏ��خjkǟ9�\��B��0�H[��g����WN\��q�\��y-���g��n�IRk��P���<�7 `�n��%>��@lw��0�����ܫv+�R6ZR�"�e_����������m8��@��z�Fv�~�\Ƃ�����t�M������W�uo�����46��a��R����e!��ɯ�y2 �� ;J�3J�W?�a�M���lt�9��XվM�}t��` c&f�Ak7�c���>� �]�2 D�a�ƌH:�%�N��e�tj���;�w��"�#>y� �l��N��/s��q?k�� ��^4���n)ފ�G]�=��Ҵ밌�@9�
S*A�>H.���P�|��0t�Q��Q*PMV#jmT2�9uqu���e0B�(������O<4��cfӴɽM:lLx]��k������y8�<��ڀP��/�i�0X6���.;���*~�]���~�^�tW�[���j1�A{�A/S?�|to��0G0���6a����i4��7����l��H�C�
�Qp��I���l���;������)y0�n8��,�<Cbb�j?�w�0�
�+�<��4�{!�Y;��圎����{h?�l���<<aG5>��,m�z�`b)�A��a!bf�D�(� Ԓ�����<���]�c����/���.���&�H��M�T�q�sN9�6��b-�Ԋ�r���i��M�8"�W#B��u���n�ŀ;ܯ�9�ߎ�����>�WS�_��&��]1���S��i(T�� "���^��/�>�e���h��r���7n)��A��:=	�2`qR�����L)7����kc������V]�*����1��"-��<&�-A�G��x��X�Dh����8h��M�r>��y��[B�������/��h��W��x�\��i,$xt�f_�R����@� �GT�>�5srIQ!W����v�Ψ�2��RC]�°1!<�X"uy��7 `#��a�њ�L QgD����$0=2̏�-�KY�o)���'��{���c��^Zk��O�H;�/?�O�.��]��mj�e�c���\܈����s�M�Fz��ٷ<����(Ec���Ԃ����g4������[^KA������}�Xx1S� �XT�QA]s�>���T����Y�%��"��&q����%�0�F���z3�vj��\������,��m����|Wl6�Aky/��(tԭ��϶ �HƁ�d�ݱ���1o��0��ICH`�=y�k��,��$N�6D� P�}u,MtW��@Oj�|[��X���C��-��:�Ā���e�k�Z�7MtQ�6�{y��ЭyD�O�e��1@�!Q}Ǘ�ou��*y�?A�ƨGy\ ����d?[1K~�$a�������4����5�y��ns��-3-� ���g�]i�|�P:
�l�|���F�I~_.����Z�w�����	��D{~���y}Fm[��ζ�*������[��Mw6��I�G��
��#�]W��jZ���'	�nWV/��L @mc-�4=��tW�h���$d�n�w�tt2*x��pm�Ua|����u��Nq�y�S#��Ҥ��T��x�|�9��A�A�C�����,���nc^��7P�=9�&{�i4��\����OW�M�*��TZ�s#Q�F��Ep�Uғ,t�y��l9ѓN��S���Md0��'�n'zҩ�0{���ع�q:^%�� v:�-R�NE���}�Uˤ�$lq���|n@|�H�o��gD��}O~��%�	��9�ȸ��G>��b�-�r_n�:�Z����� \:��:O~� �rrQ\���lY����.��2	
���?n�Ϳ�A���UF`��k>M����::~�CD������|[�� �-�$�GN����
xF�mތ������N�K���+�($|��}i,�k�J�ݘϫoPa܊Tc8�.�I��:+U���M�lտ��JH�P"l�R�vF����!�LHE���BQ^%#W��k�LZ�c��{��l��s���{�x�\�c��R���`��*1]��{�j�?y�a�+;(_v>4�-�^'�hs�����7�{��� ?��0��"�N����u��z����Y5PC5�m�蒞q*��M2����"Q[w�ؾmzԽ]��XPz��E� WГ���g-�� �ao����ow�x��&�2+b+�9Nl��h!:`\W<dE�5'�.�4�b��[ <��~R)
銆P(A=���@g�����
7�(�bN(y�e/�N������_���2~x��u��	��^���s|!�W�ھm�P�>~�OJ@ ���,��3ی��_��_���Y<Y��/�gbjK��L����EP��⍗I�Ya.��{�
G�m-g�k�ȟ��J.�H$U+tDƳ�nM\.Az�GQ�^��f�&}���N���95��&�I��I�q��^�u�vKW3�i�
��,H��Gz��*z��N�zȭiw���Y�3��� �
�[��,1�}��	F��3u��-UǢ[�%s�?�TԒ�M�
%��*8�)Ƙg1��H'�,O�Lg�������B-��'M�]���I#��b���9��l�%�BP1�SV�V�C���
+C���l�5V/���?�6���Q&�V �Uf����G��
�9�J��Ȕ�M//��q��cǰѠ�v�K�뢋��6�ˁPT�]�@�a��^�2�JØ�᩵��v�P����V|xm$��3f�����̽�0ƫ�r�����ێ�nlb��T�ޝ��F֩�_��x},���4��J5��s��g�w�Pj�̮��C��Lvڢ��6~�%�Rʋ+���L`�5��1�7�� ?	�#X�0ڳ��}�1���z�Z뉥��?�c�L�ez?���D߃i�.��L��͵��z�P���1�qy'�hh�bx�Ϳ���[�sj��w��d%Q?�^�#����Yt�Q��\��_����������>�{��J��µ���jqF �j^�����Z6��WY<�2x���i��`�����r��0��<��=4@�_�NC�2��r���yC�ZmN�yb}��>$i�6�-$�P�Sޛ���f���~Ǧ��q��XL�"2e:�cI�����c�	��וj��J��GE�Г���ODr�%��x�6N�����_'u&E?��ғ��H�"��@e�P_����,�L+�Ydf�y�L�J�����GP��"���G�,�M(g�K�]b~=	<d��c<i:�l�$-S����CU��0�d�<��EqCG� ��״:xC9�u%���
���H��I�=�3�"�t�5[	/�}�I#�	&��"4&�,�15R�b��^{��c�]�I�1�E��.�0!{6mф	��̵�����S9q�^{O��B�[��ln黮�^�������8����B��0���9m�I�
~O��w��[ �p���M��iY衚�����
Lb#�!Μ��N�����nf���
�i##Ɨ}��O��� P[S>���nzg� �#)�����*�?���0mGS��X1�TX|��i��!����5~�`���@-m���@��?�W���d�N�Dˬ@�3΂Z")%���@��	�ڧ��s}Ԙ
z��������d��&�L����Py�V
 ���)f N�7�N��"��r�)�kmz�U�-F-AP�BNY*��Y#K�IR�<�k���"e&w��wQp�_c"�4����|�� aH��BxJt'��q��/ĉ�Пֲ��!�{f�2H?��5�u]��t���=zI�=��� ���'�*���Lzϵ8���9Qc����.=%�x'n*�W���}��WGC�+�b�x��)�n��ϼ�����qN
Iۦ'^Q�0g��S&����@��N��MW@������Yā:�;p��_�X��j۔�|��f�U,�WB�"�X�^a��V�������
:�x������y��u5� C���h��2YC"�Rhv�������u��C��Z�x��`��fȐ�n*z^l��U������L��R�è�����$l�����O|���?�NT1�f��cl�3T ykf6�B`Or�Nj29ץb,&�[�~3��x�x��@��d_J?��$`9����r���`p�*:�οa���T�LN�PH�\�Og�+eeg��/l��ȟ6����W؛��q��恄@�ew�݊�������kc`<~hA9�����ƻ�N����R%P����_�`�߼/���̥������]fc�>5�-r��Q�n޺Ϋm�u��$��:G_���a�5o�r(��On�S��'�1lfV�<K>i�(���ɱA��h���]��:S�C�?��OY#]��텬C@���)�ר�*j@p��s�ur`I6C��އ5H���lbA����"_Cx���HU�}|��2�7�	$�wz�
��E^K-��o��I�2j��˟M�׳�KO�c^��J�ķ���O�����7���r��m� ���6��%��%���A#�:�h��]*��s#u��(T
\4�(U�<���Q��T}܇L� ��m������g�dp�RZ	<��;��Ծ�`�
��1�3�������u�	.-�����8�VFz��G��d�Ĭ���F�Gp���w��+dN�X�]6Xz�wސ�Ll�.����N�~f��@��zC�*zs����.��ФP� ËΑ���F��)VO#^����FpBE��:{�X-�RXU��,=%�L�;��4.s���'��ra`2�
�`��L�Uw��ɛ�
��9 swRqx�d��(��WP�FV��)S�֎=$Ew��Q�Y(��`.�":P�����8���+����%/YW�T�#�&��a&>TGg�3�� �-�
�~V�5~i�<�i-q�у�}�qB�=�Tp_�%��`\�Ffءg�X�]t�='�H�C*\J)���cXu�$!�h]Y���z���U�~�<a��!RÞ/L�_!\M�4d���S���e��g=��!TVqߤk���T��\ՠ�2�i�^��<��O�ʛ��?� h7�w��͚-���>���'��S@��o�#~�;NӰ��K��x������6�Cv�	���R���j�-J���鑃o�-�G�%�*�N���.����hnB�m�b&�]gw~WO��T�-�y3��Q���&^ş1��X�i%�;੆�>�P�\qn%~�id�G�y�`��ۇ�t�4������[}�n� ��d��-�i���h�X�w�W�"y&˾P���B�Éܫ���N#D�Q�o>0�q堫��G^$8�\cLC���]0��-�"n�(u&�=�{� �{2�ڡ��gr5?��;�'�P�8L�ɰD�#sμe����%�gQ0%ȼzx��wp�b���/��&X���L��]%J��%�g����H��i�
����)�>&n&����@K�"��i~1�����
|�><٧\��Q�=���Dy�~��AC�6���=�	�$��F��Ʋ�W�Şp����%�&�:x����K��9�W�ZRL��FVsҌ������5���r@����ïH0�A��p��Hw�'uP��_�J�� +�>`)��!1�IF r�O>E�6=(�#��:�r9J_p�TX�HF�t\ְ����R���<�:6�1��ׄ*Ȓ!&��D��?��m%�����K>\f;�ՖO���W��p7!6da����@��Q��˻�Q[XUy�9��xk�\+�N?y�ڟ1n)[�c���R��P{M?�dDm��pr���c����Ǭ��%{r�B�b'oNBq[Hf��b�(a^5�
T��0-���&��hg���Ś��w5uk�Q=f��� ���q��c��輍?��*S{�n�x��J��$���Ś�SqY�3���85�EU^(W��-��+߻���L����Y_u0:&�]������pw3n�,f�����횱n%9`�e3jn�7`�	���l5�D���+L��?�����|V�����ŢF�C�2� �!�
�����w�TN�I�K�!i-�x�a�E>'� =uV`�VOOM^撬��# ��J�q��)Z�2���7��́������p@?69^'�e��bF<��b�X��\�UO�c}�8f�ڈ��_D�����.��}���?��8����Y�������Z�Ue�Y�ݤ���b/5m5�2`��]�	�O���)@6�;�s9�@y]�@j�i��YdV�D����\C[��?�_d�� ;,�`*e��0����'e��A�)1W�[f�!Դh��K������,d QѾ��U>��5pA`75�o�4oS�p�ؤ��A[ó�0΂>~3�{���h40:A�w^�"%���q0[�L��F��*ž��S�p����
�Q\����}W���|�@��b4�ҍE���B9��"q  f�k%�\�'i�����D���ή�Z�����Qt��j������m�W�\vS@#���X>(F�r*΅����N�dj����|��>����8
��@Cq5�uG�E.:�<����wBs�� �|�P��ҥ�Q1�퍎U��?�I����%��=Z����RE�p�uφ
�OFByKd��5ɧ�(�$�X��Ǽ��8��	���N�,�pD�D"���e���}K+z�{<�j�|��qIz����E��d��\����ʯ*��R��/�gck;""K�4f]��1��X��	l��cN�_�}<I��?^6.���,W��iE�	x�*�Ҝ+�l�x��j�8p�3��5��sr��'�3gNs��^H� �v��o�rn�b6����·i.ٙz�}������`Ec�x`T�/kd�h���A��ME=[���#�NՒ�����QR������~�֘�c��o�2�	w�vE@ւॿ~�m�[-�z�\:��#gb�b��8P���Q���7G�.�,��¤�n(�����߅~�5^���fY0�2QSHa�Z0��ԫ��S�G��}�UIfޡCω�ұ\@�����ѓ��C� f�TO
�L�n)[r,�G��q��jw����V<��%n���{j��'�k`s�Q;�l��$������T8g�w����|J��8;�?P_1B�6�|�Vbص�����2	1�sA�����
y;� j�)|�,&U=-�ITb5�R��s��\��\�?�nP{�9���$؝���#��p���^����.��w���2�k�<�B	�0|�}�P�z�FO¦�B�AβrE
=KDRe�1��%�/{�����.4G��� �{bZ���������TPMɵ�V�;�Ih}IQ���f��~eJ��zp��h����y��]8��z�j�j-��&�b���9���8��jy�d���yF[֤O���@�#q��&�8����TZ���<dE��ˆ���_ʦ^�p�ǭ"gF|�ޔ;�P\��[�r���9D�&�b����(�Ysy��t�bQ����o^
߷F���5�E�;G�C�q���y鲐@2r@��U�Uz��wEC��ڹĆ���[�[�ZZ9;�C�Y�)d��yd�&�M�G#{ #	�i�$m��C� �m�3r�Ԍ~�i�ó��홍�8�)D	k�~��	d��l���j�R�����f0����pu��;������ hT��D��������/��LS�'cE��}�ݎ��	��Cߊv��h���r��" ��X��+�r�m��Et"��}Ǆ#��m��c	K"����sC,��� ����h�iiIj�t���|��\w^��\����b�ٽ�żԜdٮ�0@���59KU���]���ܳ1�'�T���8��WB�Yo/���癊/8 <d,�V"'#��=�Һ:��k�(-���ϐ�ª/*��G��B7K��eL��am���:���F�X�GKJ�k��� 9��3'!��<
���ߧ)�X�܉�)�������Ei����$.r�j��R�1����J�t��}�� �vt�gK{����)�-@���S6]��G��ˉ�"O���E���z �2��X�m�t4��8�����a�T�~��$z�ܮ���E����� �xu�N,,�_W��Jn�>Z��2G�F�-�9�pm	RP)&�xN�T���t�� �Pq�����(�p0��t��Tk��!��/=�C��?���Y���q񱟇��7�Yܙ�+1�؋����TJf�#�#��j�bĄb(��4��-��ʨ���p�(Ǘ�_]��K^1��_A@�O�wybin��]�7�9���	=��6���0eg���O�<�D8�,��	9?���
KQ���	��i�YZA�ieP�.s6Xk	F*m-��Ձ�.J3E��sY����@1�2�^��?lFJ5�)#�'&�k�-���TǡF5sJ�{�q7��ᏚS�.�ٝ'~����S�ha���w�F��b���L�п�d�v*�D���G�m���_'Y�`����(���tvqby��1�7��!�3��}}�#$���q?�F+�Zi�f�cl��=��v[��A0���wL$�1�I��w]�Kd3Jnj��Il�+ã���`f�9�Q䞔��z:�����,`T[��:��_�y/������T(�7Z��^��a��(�X��xK^��O��5^��$�}�Et n�޺~P��ۈ�Z$OŒ�&p�ƥz
��1\���͢~9ڴ�p���#`L�YJ�=�N6�N�-�mY��Q��5����+����d�J�� Z�f~�����3�:���(���*�t䵉4�uC��w�B��#�����A��VhPt4,�w�X>��Vʬ� ivNC�X���o�b��Ӛ ��a!9c٬�de���.��vN�UY8UG�����j��g�]��Kn���~
����x��K��z3}M�Z��aQ85D��a���@���5e/x5;WV�	U�O���G7M��FO�U�š:ʠ䡄S�\֥K���u;���[/Q�Ё�t���W�#�8�07Q�	Kٗr ��:�n���ݣYr�����r���<����7U��ŉ7����RNC��.D��n5���]��/D���zPV�˨�!upZ���RP6�+�~i%��k[�0��|r'\u  6���뇓���n~�S��]c���W�n$�8��`?�<��ܮ$�+���� ��N�1�>�OG��R~zYsľ$_"��Y�kh�%��V��_�3_��\�G��s�!�X���M��r)�%�l�����Tۼ��_�[Au��+��e�%0ݡ�jn�s$�c�0TO�!�Gu'� ��juɖER����s���P���~W�9ZW'Y�@�]0?q����M������5{�ޞx�k[X9����_iͶ�O���Y�� CQ���8�	 �R^q[ͧ��1��*܀E�8������:�U��"�Bݼ],�zD9�Fn��Dm��7tk2��n��}�&��|z�
��B<���ƽ����fV4|�a�.��:�3��:�
�~�1�(��#ǁg���OabT�.�ꜻor�� �_��;���Ŝ��G�J"w�$�	�'�������~ж�%qyR����>>�|h���J��DL]��gR>��)�7ƐC������lp��3S��s|fϒ��Jm�ј�
n	�8I��h�1NFbJ�.x(B[�s����3���j;R"wˁß���^'� �4�����>������P>�d���T�T���$��� �,@ԦU]�#���37OL��ܑL�-%+�Z��풊KpuL�]��*lky��
�I3<�?�6���y�t�\ �/4v.M���׹��
����fr9cF��N��b2�@1z��~H�l\�?�4� I��N��� uV��߅�/�q�,����0�v����u-����Z]�6��+���Am��ϡ���X���L�����^IRT���r*{��a���3x��k��p9zf�r���1����¯np& Y��=[�����d�����?\�+o�U�L0�7n��
BY'���rU۱@<}`2hV��Sd� �X����fP��Ss�e4іS�҅&��9�i��p������?`���O�6v֧
ކ�����rv7Q&A�J�w~�&8JO_������ ^�@���H�)�̧?{)���Ӎ�~�1by���R�	��G{	.l�MI��_����V��Ud}�G(���"�Ԩ����R-�Zٓ�Ѥ�p� B�C'֠��褵�>;U��a-��d�B�/��7�μ��F-���<q�	!�Q�Y-��f���ه6�� #c2'P�V~�|t�ϒ�,�ҳ�Q;R��g��L�Wm]��V��������Jk[%P��i	�E� ����Tyx�6�gJ�xa���� f/��!t��~<��KW{���2��М�� uz�U�45���3�ڬ���Vu�IHMw3��ך⛎C�8� �:Xy�����Ӳ��cLT�K|#9gKG�e$qj��]{�9�z������O��V���ߴ%�\/2Ğ��<�A��}��������Ju� H�cS믯���0����P����=Q!���"R���ş�L#��~�(�;�%mHs��*�g���t��-�fb9�+"��h�sj2�g�ߙ�
f��&x�)U���N�_������}� �M��&�cS#F_��5-�cfpM8�?xg�i�6�O����}l?�����	�l��&Q�QUy&�"%�Ff��2X�!�����6���!�T.���OC�D-�`)m��z)9�!͂=}`�O���La��̓1(ZN�󯗾_d��܄oR(�B2L���^A�i���r�`2i������)" �gY�k��(/e�/�������s٪���w��mc6�d��j�(��l�+��5=����3_�^]����Gc��`*7c�7�Ε׭��4������y^f���=X�����C
.���U�KƓ���
�.I��-��׹�)�d��6��_����]/)L���4zn\�LDf�����z@Ǽ���2f9=�G�&,�a���S�6(�c��\*�Y������)��0De�L���3a��g��a�.�.����F(�
>�9�Bx9f�^KPHl�	i`h��i�Z���h���� F]���F#1�M21)6�c�S���yr�{j|�7�+¢��Z!�5g�Ҙ�2F{2�Xr]��H����05����)����U�	����^��k�]w'�{����eo��YC��	�=�a\j��_Ӗ�gP9ޝ����t$��g:8��#z�%z"'OT��e��� /�[�$�ڂc�7�Y �qj�l�ŒuV�/�W�0��E���a� ^�뀡��+�74��{i�W��n��LQ���ހܷr�>̾i�˙����V��%:���Le��p�ȃ}I?F���v����+؍�Ԥ;K��z͊Cs�O�5
�m����Y�IJX�Y�5�(踂�(�s��|-��@K��~Q�Ѵ��=��!]�$AKzH�^�뺲�{�2��8��c�n!�z�w2A��06�H�8�!�3Ê�4&ya~EX���\�r�JS�gn�J��]x�����K'u�����9�%���}��y=�p��_N7�V��׉��P��d��
!����Iݎ�Q2�1C�`�q5X�8;Bq�ˮ�KE�%��{x��8>Rw_��k�8��K�>0��)�c�䥃 u��|��|Y#���s<�'HB�A0�O	�������e.��")��Om�5�Qw����`OT@]����x���v�� ]md~�Fo��/A��I�Cr������'B�==�5ҭ��b q+0T���B�+�8���	PR�&�:7v�2^���N�;�(�ڣ�r���Ϧ Z-VZUus3U���%C2�r�p{��ůX�23L�*�g������1�.#m8+��M>���d��caJ�I���FX�V��cB�P���n�n�Bs���O�&�P�� �s)�MU���X�TUg�%��4���Ȣ��N�X����&Vs_��	c�M���EX�	�+.�t)�Z3��h���?���'�-�kx	7� ?�h���6���7�>~����n��:�9`��C���T�}�Z�����Gඟ��� �Vꦬ�vn{�����b�d~����FMB���y��&��N��Y]~��.Pg�M�a1){������م���Q�#i�K�"���J��"y�1�g!�s����5�ғ�~d���}�H�;�'��J/�c��(&i�1��IBR�Ǎ,��#���7�R�~QZ����f��K�6|�{RC�� f���� �Q����Z\�P��ܨ^A�'* ���|�ߓ�-o'!���_��I�C���a(�B0U�ѓ�l��g�`Yb�m_2���p_	6��v������W3�*K<=�7g�KFi)��@$�8D2�����@�x��g˞WA �u}�=�8�x��IR$�)�I��Ԗe/��1_V��e�"؅A0��Vݖ�BD�\ң�*O��1�d��_:�P����֎Ŀ�GK/գ�Tf��i�N� ��MH��L�����Ie��������c+�U��wn�X��Q̋�W4��0���h���h�(H4��QL�R���5|m�w��p1*�R׶�3 �s=~t�6�w.�$ScJ�;V���o�q�8p��,
Lo�mKP�-�fr�S���p瑸%�~����h9�}O���)t���d?��ڥ�i���\;�
����N�����Z=Y�OQ�kی�̚/V���;RxݴPX�x���1��6�	j�ݿ;ǘT��U��% 08]���.~��E��Rd���PQ�I�v�9F��f)%��a�{��I>��6���9UY��d��f���w�7�̀gO=�{j�q��ЫA��U��Кid�ZH$�/���HI�o�#$�K���پ�B����X�H��!�u��F
�ee�EK'��G��t)
N;�z2��r�,���*�&�#��v ��^,��q�������I�O\Qg�+g��i�%�q��n�t�6j��d.�e���%�@7�dK�9/N�}����FjH���*�p�Ui�g��C���o���u���*�b|�.�`k�Gg��. ut%��,>pe�O�!Qf,�D��6�-.���d��z15��J&�g��t�Ⱦ��!@�������<;���ⰦPm6e��v��p�%�>S�� ��@�G;�D2�P�\��U�~�-�Gp�j=���Ox�~
䄜c;���3�������N�Ł�������jOVрi�$PB��69�}��R���]u��8<�GF��I�RV(Sg1��]�no$H�ށ����vX���3�ě�����q�Q��^ӻ�+)�@�x�nEU�(�kZ��7S
���^��Q�.Q�bՄ�d$����SChqt[����o�Yt��[���,���뾫R��5��昼I�r��$����Y�t)<�n�`w��Qh��PF)Q�k�.a ������<�C|�+e�R�Yy�4�i~���8��4Nۙ�N�+"g�J	�2�\�6�6͟qx��j;�iqU��{����GWhr��U�v��4��i�zNۂ��M!y.��]�,֜�<�%Ӟ�2��ߴ)cyզ�`T�-:a�K��2��D��%f��%�%Ys�$|��@M�+��I1����P�����so�0���yf�Y�Ee�/>p�
��F���("��u	NΑJ�:t����m������ע˔*)H��Z�~0|]e�)�+�K�I<��6-���BH�J$g�*����/O���<#���/^ߦ�8�����H�Ҏf-M٪۩w�`ӰF����u�ψ�{Q����:N��C)�������iu�,�dݓټ��B�Y��k�A�<*�\y�]W�\��+`����<�$�Nf�	��Z}h�^LVڃ�nH���t��u{��=j�8�cIe�� �D���n��;���#�:i[/���$�?#���T��U��Le������.�I�?c��)F�n���c� �T�"򼉜=�Oi��"���x~{Y���w׏���l̽�|UVAm�n<�d>��K,$P�W��a�'I�}�'�w�m؅×���:E�d=Hi�6]�8I����jGPv�u����ߑ���'��ԭ��f*>�tb5�f��Y\:�oW8o-�ŷG{�RAPL��(9?{���������s��k�ˑ;^�$c~�;����=թ_�u<�?ԍr��e��c	|\�%��Z֗ѥ{�~�q��%��f��jC��m��]�Dn& sa������h_��
�?ʋ�V���~���P� ��T��9�MX�>aw���]S�y��r0�h�nt
Q�\l*�V���S�e�aL�d��~&�+�}:�A����d�f��ŗ;*e��sg�L8�ޫnt=���[�O�*�瀃c���Y�!"�wK3�E�Jԗ�P�Q�î�J{\r��O'liN&�5.tj��z�۫n����~G�����'�|�6W���ؽ���]����h\F�D_�J��k�ć�9+)�{�	�dTP��%���1u8�t��Us�$u��)|��l�5`jF��xnV���8���J�n���M֙�\����T%p���uݵ�)e������cv��+
���TR�?�)B�L�o��<Y��`�����	�2��M����.q�0�;t=� ��p|�� ��nm���T gW�Y/�Ƞ5��1˥��L9�>��Uy%2{�J�C�tA���+�q�>F��ˎ���H�PKW=[����,H=f٢#vÉ\�ki��)4��f�Tߑ,:���æ�+�Hd�͇������Oq��ᔀ����U��{)gQ,?�-s��u�'��2��N�3��x�h}�y����k�I!=aqB���A��\��ԁ�Ӗ���v��Kb��P'?��&r�M^ل�t�"����t�2
�4��CX�P���fw~�N� J���"2ߒ���>�9��S��y	� M��U)�H5�匶��Y���gH+s�.Pz����ֻ��_��O,�f��,k8�.?�`�.���CS��ɻ{B1�	Y�����H���Η�Q���U��lȲ����W,�v"״�J��d����\�"q#����n�퓆G��|���N>�:$+�
X���mε慈syXw.���"��lG���A,zD�Pi�J��#�(�ߝ���Vڨ7��#w�ZrX��׬���X�`n1�x������}����՘�X������=�:G��wQ���4�/���!�х ���u����p/��ҁ�(XĂ��"ϫ�?f�>/����3.)�AR-D��Q]t�.e[�1����Ûd0H��Y�+��l�tgmel��
�=5�L�0��hT��ߜ|���/]��%��u۳���%����5�h3���>L�V}�/ϳa��:��{S�c��*[�
Ѫ�Ae�SO&q��;�>��Û,	��R�
g��g�*v-y�71~i��6!��{��F|+��*���4���v�ڋ�g7��rN�r��$�Յ8�( .��b��!��@7��nE)o��P]�)�OCD�{�#����vm��aځ%�A�2s������~��	���W�UQ3Zs�"f�)6�/+������k�-Lw/�Lˬ��_P����DVB
 ��pʿ�?�� ��v�y����V�L �6X��|�p,עr>�.�ʹ �Ư��a��2�����x{�R)'��y4��{���k9 ��8*��^+��O�6�DO�ș��7bs��YKX ;=~�U�S��c�u��8�Ts��k��;B��B����ˍ�nj���*�@	%������WZZ�=	�v8qn�	ы!gPLu����i��C���",��`=D�,�3!,n�\���<��j=o�w".�mX뉘$dY��C{De�LB'�K����87��Q�"\#0�(vĂ���PK ���D�Ȯ�Z=����>[8�ӠM����m����7xTvC�8�W���a+�@.h�
j�&ǩ�����m����-�2@k9ŵ0�~�,"53!�î���	f��t��R��G&��ƛ5�����e�:E�[�G�%�v��KFf���$��K��A:g��4��%UL��B^��T��,oC.�]T�/~�~;ܥvxLP`⣫��t����&��������5F����8Σ�G��7�x�9Ӹ�)}	�P\�Kgۗk%�M<����z���[y�.������!/�V����"t�.T��E���w I���v��P����]?|�"�ģ��e��k�A�eZy%Q r�Vu��<m+?ɨ9��!\�Z��їR����D	�~{��`6rYq�6��=�߉r���b�NBT[��\��s�����?��bi�����*v!�����b�P������#UL��v�a��}M�E?^�P��iE�녛\��Y���C(��ï� �i3��/9&`�V�1�N��S�ædu�����S&4Z[ѱ���'�Ǵl�Gw�=���^b�t��$��p!J�ѩ|eD���qW�s���)�|&�t��|h΁�2~�Nz�-�����by�S~nT���I��֧[��+����v����jUM�jx��Z�S�.E!.�7�����![�p<|�9�)^&u�z�
�ӝ��h�����7�اa��n����%s�Rƙi�$��]SM�@����̫_�^����(�4���_?�$L�SOy����� �߇w��#��J�	�E��%���Tw9f��J��t�e~h�u��P��#��tm鶒E[�����V;]�OZ�*K[��԰��\4�|��?����Z3ٕShtʷY�Â�����6��%��<j���H`RUb����ZN���#ڌ��W�i�e7z0v�=�q����Kժ��X 8��N�O`�i�*�6żS$��oO}�%�OE~�O������HK�kצ������|+-k� ��1M��",B�{�.)�be�C�HE��m�5^"�`?���n`��p����N�F9'
�b8n	������xID �������ڋ�л9������@��ڭ4h=]��tmf$��#��p�3Eє������!+@��H��i U��#�m*��:r��y��rMJ��9㷗q/��9;���j딳v�̟��� ��Q��°hPw�ᘐ�!t �����v�tIC0���O�lm���v+�:�sC%i�ry�K����@b��y����YG
p[Zا�@�iVGŵ5:(���rY�hh�j�E�/G�x��oj)�I�D%\��U��H6���j���7�#=�.�qp%l�W���^+ؗ9�M��s��Y�+}�(ު����J�}lw�|���r�4��VR�����qǱF�t�iYx<kFF6���6�^��]��la` ��j��b��"bȼ�Xv����+m[�z���1��D�*��������ew!)��r�W�6<��Mʣ��=����R����Wv	���'/�(kR%Ѵ6�X�hE��0����8y�bt������ر_My��D�/�;/��qX���xʪY�X�V�T���ӄ�S����v��=Ԙ��ٶ{#�A4|�~�x�&i�Q�ŲWP
��������.��_IPba�:�?sAj��M	lKdV��}�� �?��,�9޲���9a>lKP%�BòW�I~R�B<�6{Z�k�uK}��*���0֢j�����\��C���`�j_����46�رn�]XY�_h�h
A�+m�5�Q�*p��5���,��H�dG.�����*
"�G��IsR)�q���\Lv�2�������م���$2c��Z�yᬞt@� W���
E�t�f�g�z�e������A���o߉z�独:C�� E�*�猲˵�-�o��*K;f�.�Z�H��^�뤀�L�y�$_v�S7�p��#��Y$���.|�Aن^���L0���V��x!�>��V�j�����Aq��xwM�c��{��� c��֢Sdm?�^��K|�~x(�U��H��"c�ʫ]%�5�\�_���h�}�w���A��D� B�ĉ�����@�s��NjI�y�Ј�Sb5-��D3��GL����d �zA���~�i5mt�"�)~�.jP�٧(�:3�žΆ��WǗ��"ª3:���}^��e�o]D~�'�|�b/]��=a���l�N�B�uoY�Bɤ?����a�<�/J��-7�f+
kp�E�1��"��[�^��s�r�g��
�˚���Q�C�����A�F���N�
�wDK$ �E���:FNE����^)c�B��.���>���}š�fu��>��t�{��_ͨ���Ȩ}�ȋNa%�M�Bf�cv�{]�&����j�?��N)jE��HV+�W�DL�h��%����}u?��"���M��?`#���%��(�ZT�J��@C��P�"m>�%զ��$v^�sZ���Dv����}��E��1���k�5�~r2���,�逐fB񪘓���'��5���3ef����C��ϴ�������0��Q�-�ٕE�۰���A��ˇ�f�eh$gp��nW,A�K� ��hPi�K����i�!=�*��?�"q�k(?����E"�.���2/�'7�-z��AdΨ�G�Rs�)O0��`"��	�N�$�-ⷈH�Qo
{�[��7q�V�����?u�ՉI�3��v��8w�0�;���j`� �%Ɓ^K���5�'N?�"> 'J��FҚ5���}I:~���=�>�����leH�D=^Y��F�: �8:rjr�HdV�%Od�O�����˄����WEG��d��[N(�6����F]M �TG��UPh�0�$�����o�Z��/2��"�ݽk�AAP6���9�=g��imu
3]�;עd*�@�G�S�д�Y;�� �t�=���c<����c��"�w;Am���f���4(��.���<.bYO���*o�m�0��oJ�yXU^#ZE"�3�z�%�&�d��#Q����tp��]���S��1^�ӌ����b�''&06+�����x/; '�����WO��d���:+�d�KB��Jܳ�_�!Z[	,�/��֮]���[[���h�v�{��;�ݮ�/H�w��4��k���Q�Lܨ�]��W �cy����__hP��5>�?�BxC�H�'p��^�Ɓ��k� sS��ﱵ�`�yy��/�?js͉ �E$dR��T�3� -���b(�h�mr��5#��x���լ�F��a/�����#�q���i�vP��
42�ځ�����"�Y��'�ܜq�+�κ��/�Sml�w I�s >ne���q�]O*#���_�R��N��]���-=���d@��0�Q�qq�3�:��C�wr��WBy �P쑞!�Z���`�јV⻾*���{p�]uةk�M�����cpJ�Hsg���+��%]��I����_�\�\�g��E�����g���=�~���%p.ߚSf�]M��d�~`�TUS �;���7엤�1���!��L$ZA�ts�@]O��	9���j�U^e?����v�<�	Ϡ�{�`g%�E��A�%�I�-�)G+*���EB2^Ґ�;�WT����`i���a��v��<C+V���^������Fۻ`�p#:
&�њPX�V�Z�0�$���}�~ �^~�Lx��"�u�hcȸ�^�x{������3�G�dy3������P[��+z��Xd�D�U�Kh����q�Ύu+ǉ�#%����Fƈ�~���6����K��G��2`f<�G�h�4�����ȯ��HpƩ=��3h<���SE�aJϏI-�x�
Jk@E
�>͂#b�urYP��
`Ur��ôFk�B��ÿ?�>5J�w�� `��L�֚�����6�b�$�{�+� ��u��X�d�9^�0{��;0
m(J�E"�_��<�����\�D��	$�.ϷS�~�탗�����(0|Ŏ��_��Z|Ѓ�������U1eDN.��T3[k�����}���:�"�"\�I��,u{\օ*U&^��Rd�:]�!�Ga�� ���"����F��ώ���{��h�쭥��%�@������CP�I��5"ۮe���D��W$��b����t���lx���'���̘`���K�Xg;�� X�bL�-ED�[�t1��ȀYr�h}\,Q�r/a�z&ecNA�'��2j-�w6鴬@�g���h9�A����e/�˴��d��s����NZ"����`�&�ZI�m�nU����S�/f׫�O0�B^����\�y��N��>a����"v*���[f>���+M"�K�$ACW��i��F.�����?��6��Zw�����B�rW���_��m3:�*��1}�T��R������	K�D�8�m�BjJ�ti��fb��Z�f3)�[c��M���o��]ِ�Ҿ\�!G����������]|���]��l� �C+FF>}B���g��S�y�H����������o���f;��vW�6��q�ݰz�Qa�Ґ��|�%��=x}2���5����ٻ�к�l(������.�'�;�_o�
�7���.&T�.�O,CCR�@B
+t��82 $_��1�C�1���GAn�2�t���cB��k�/Z�����ƣ9�0Y�
���M ��sr�/����퍳_���>7k2�	�C� S9B#@_�1{X����1B���J�וg��ڃ�h%u��\���o_X��h����A?��?e��Cj:Ñu����Z�� ���e8����u����Z&=v6CΪ��l
�zc& �?�n�����8TrU���dp�_��+�E�:)NUC�D\@���
P����\���e�	�#�8�҆c�ϝ%�Ug��)�w��D$P�zw]9��{��c*簣�b҅Eqo$�+������r���7ׂ�i�4���|�ۡW��eԤ�3�lX�����VO(���T�Q6�2�R&|����Z��mӗ,�zd���AI�u�Pv�ϕw�T�ׄm]��T-%K�����ope9C(*+�VU����T߂/��|�'�Ϻ�u� �zf�h7�����Ѻ�(���2AK�g�_��7H8�4B�"�y�ǌ�m�)��E�Sz%�uTȸ�����.Ipnn`/K;9�n\귿)D���	�D,�Ӗ�$ƭ	Mzj����� ��&{�KX���$rD�;����H�k(�3��!K���e1��>cv��f� ���j0ta^�8���,�a����&	�|#�����Ϸ�?�'�0�$����'�)�D���4j�ݥX�]��‏v��� /uV���_ow?hD�Y�$��(���.ຆlv]�<�l�n��;����������G���j��~険�L�w?$�g:Łzc���HӦ��f�Dn3�u
5�u�Ly��'m��Q`\U��J8���&���N�3�*�r�1���>�H��T.V�[x(�tI�>%����p���f�B�m$�jT��P���3�~���eS�/ 3�)K�O���=ê+�W�B�,)�.�h����A��V��k�Ҋ_)�;Q�E�5�?-����n��{�Z#�	d�	P���>���M�����@/��&��	�h����0��ٰl�#Mň>|S2��`�W�U[I�"F?V�N���~z�4�말�����J!�q�]1�H�����N	_�f�ǿ��Rا%G�Y9K��P��^��ju���YR���HV�&�Lp>=��)�Bt��談��Q�yBM	C矔�[7$�+Q�1>�����[�p�pVy��C����}�>y2	ұ@g�I��*\�u���W ���ʆn)6]P�c�Qz�LN��fҀ^G� �&Ӈ�DR9�������ȓpZ�� #?�V�mI��@#l��&��m(�Gcn��K:f�/�%���d�6F8�vLP�����UN����/��i��p���"��v�����>B	:&Y/욊�L��IC�Z�y��vǿ�<)](.m^Jn8���3�k�j܆�,o��|Ԓ����88�gȇI�h���l�[A�ElȢ���n1b����d3�q+P��8��E	��Z�X!"���i1#�g1Y�.�w�G�pU�U��	Z5e��6b_�y��cw���!��8��:�RZ(���i���6q���>8���5tN�{n�Q�g�?�=7V^ ���p]b��g�ЛK+�i@k�Ю���ʅE���?�����z�?�e�YEb�'X}���� �����s�U)��u	t��oj��xL��PgQ�.�.�[�u��B�ǇPO/��4bby�֍�4��RRM8xO�~�U��U�l���.���N_�M�yri�5���B̙��[�$��(pVp~��E�_he��������x�o�gdDhQ:}Ɏ�bJ�#륽��"je�`�,����+�MF�ҙ�#-�9�)�l|�ݜɮ/��\A����#�����@M��f�҅ij����<�Ư�����w���{:bd?� ���lW_��$&�`�g(R���DǟM�%��T�ϻ����<&~%�"oC�aA��']����!����a�q-���
�F�
nYY�)�iÉ��V�*'�?<9�0��}#�Eی�2@w�����Ԇ�wvE�����b�l�ś�>�n/�з�g(�(���+�8T�_��7қ���	��%�[�}�͟򐺨��'���"���/�@}"��Kz{�Dɣ�Nfr�F����t<j���$\-���ұA� D���3%��r�{���M��-��y,֔�C�l'�D�/�Q���R0����͙��>�7��Y�����X&�,P�w��M,菁��%�K��v��0��=��>����-j"�Ԣ�'O`�����r���ݔ���K]X"M�E3�)�hd{�0�p�!t��0Rb- lEF����]G�n�j�"�3�u���h�>�����G���;��k�D#5R��l����N��vL��nh�!bJ����jȸ��5��&�S{y<��1m��m�&��cT�췤K䲂|3�}�A�L����<տgʥ4�������M��*{�.�I1�I��l�l$B�P�݁��oF��[3؄hyn(%S�?�����9k�`�r��T��΁tC��͘��f[]���IV�o�I�0H�e�T'��$Fn"'�,gK��Iq��m�YO ��!O�e):��=P�|�8�����2�7��^��i�4���wc��?ԗ���!�c�N��ѨC�xwN����Z$z:���zh�!��h��8յ���Q317C�J���ka�����T�G;!ߺG���Y<wJ�����0���*�ƚ@�p�F4Ȑ��m�G&'r���&���^���E�BV�7m����b�Y��%�L�Q���%=��k�Hm�Z���W��jO�����-X��vx>���]�����HLfY�qfxu��\=J�|���Et�|���m<9��G��e�"$$H��#�����������C�}|N.�$RP�����ٙ����$a����ё���[�H>1��v�/ͤ�]L����)dJzt5a�A@T�!�҅�Ԛ,6wp!�i���^�P�C�A^�{��F�=�~F��M[G���ɐ�A��	������p�9)��'�i>,�R׺A&A���s�儑�n|�/��|}u8���n�501�`��0^�hJpb.B�/��r�f�Fޣ�<��<c�Κ9���fh��]cd�2构���d�6� t�k�?ie;���g�R=��9.y�~�=�O���	!s���PO˴���=ߥx�D��+�w?�~���Ei�l�c} 	�i��9��I���/	����y��*@�WD�k&�D\���g�`:ˤ��1���X�B?�hD����������Ap�=�UE�Q)o���NWf���6�e�lP��Ri�l�ت	��+�~e�-���h6�	B�/wc�M%�K^8+m��Y�ɫت��H��;0����A����4�FW!V-�NR�=�i>�D�8����uQz���4gm!�k�j�Lo�U�#��\�S]��s�/9C�	�ja{m
���������=**�� 7<g�ĭ��VB�6�J��Cd��旊����EL�@���ÃQuQ��QK��b��<m+7W�J�	T�{���m�f�����6�CC�&���0U܎�U!ғ�������>�]uF��N_;�G�C_�?>.�p���r�5���*�X��k�[A)�0s�;>tZ�RO���D&������%�w�-�5%:�*7g�s���2�в��8�x�9��<������9�9��dZ�p�wU������"�|^��YI:����>���闟zK�����*�ԫ�����#�ڠ��K���_���W6?E�h���_d�~Q{��Rvl��&�yh[�%s���|:5�[M3�X�ХoDћ���?�-S@w���<��^M��+���ge3��h�[Σo	+M1M��GJ��~HqK�DW5PV�Z��&�g,��$wu��� 4c-Jm�Q�m����EBlN�0�ȵ7��q�W=��N~`�k���A��l���yC�`ԥ�:%��^S\VK�.�a���`��*�ٟC��NG�����(*s�#ev�s1�~^Ĉ*A'e�vk!��X��D�_�]�����b_b*�;���#���2�ؖ4&0��|2;A����yuk��j1��~ �S4�)2�[�Q*K����+�N{ s�-+}yeN?��������oޖg����pw���i^��h�N�$�d��/�AJf����v^�N�[�m��)�7*QP��w�Xf�ɶ(��vKQ�F�+��$�7{���?[Y3�[r�o��1I?��a��b�=U["��{�ad�^�C���@�,"K��}-A��]�˟O����l�f3�ɻ�h�vs���H�$���Y�L1Sj\�Ū��9���Sآ�,O�:��>Z�v��w}��C���=.��q�G��[�&m�K?�y���n|�V\k���Q�F�>�J�Vm~���/��a����;�HYk�j+`��A�eo"��I�(�g�}Xm=:l�p�/������eN�Ȕ��y�R$We���G�-Ǟ:j�dҕ�����W�}me�K{eg�SNr�ґ) ~x�����c�Ub�K�ͣ�ܦTp�88��#}
�Jі�z��/��[�Y�Q�Ba5��k>�1�	��ca���b�hLL���Wt�ެ��YI'�ߴd�	�=�`��츿���p�����z�{���߿�u��4'ޯ��_���(e��c�F?r�X�X�ˢbդyŴ6��@h<����>���;�yDX|��+V��c�ML���~�
 30���H)

�g<��~W�$����2Ǌ�)�6�Ж����4X�G��[;��#F\��/fF��+!�����r⮠NmoE'[D�J���E�OT2;�E�5	�sd�U|䞕Ƨ��6VQ�cFސ9Z,�Ƹ���g���m�R7��W4\J?E�xɿB����[�3��C9.���F�>��1��[��~݃�E�E����B��/�c[HͯcK�.�R|���w\��\a歨g�˄�ic���x��z�d6jX����kD�'�zƵ��S�B������1R��@M�z'D�I 1��<}�6$�;��]V�����o3��k)����SA}��ZEa\uFP�L(r�
�7��/��c1<��@��N�5]ބ�x��B�)�wZ��瑃��x�&>�q��]���.�����b�@�X�W&E��YG��9��gA�e$�H֡-t�9c�JZQ];�~�O"-���]݃��D׮*�ޘ߮e�ݮ�����[��o���R�����"��W�7 J�E������� #�UA�=�����&���+����e���i按�0��������@^z}��y9���m�C�`pP$����GU�:A!?�òc�a>I�K1Ҽ����
�
��?�`Y�_��5N�ċ8�>�ի�]`�6XĎ�]�e�R�F4�������߯�ܮ�^��o���ri���p�E��p1��\��=Wc��e�p̲ô��I/���w�9CY^W��z��y�Ҩ �H�t���qcQ^O�1
��^8������ ���G�&�[g�[�����]�8��H�ݮ�2�{�S��j\@�$[�h��2�\�~vx5␶N8��h'�^�&;[�m9(I�\�|
��z�bF*�Y���ԛ<2U�H�ٺ/]?�M_>�ˣ�]��p�wÏJ.�l᫋�dSS�w�2�+Z�֙w��Ji�P�}��S�M�j�~T#(h��� ��>��	������t��Lx�� �S�:�F�ىGH��3��UdHأ^���	����A����&��w2@AP��iPmr�>6�.�y���뵓�-s@'�D%���F���H�'�DJ��u�;V��&`0�(�Fb��=%���9G|���-�N����X�� �)�6���u}�ie�<å�g�B���'L�_~اR��g��O��r� T�B�����a���+ $Kϩ���L�]-����|.���@}R�3�|��	߲�y�V
f����[��h�Q��=B��n����Y���U�l���<�';�"�Xn���q.��`,�u�:�X�I���b���%�u�.WA+4�?���b���qΈ���{6.of��1�h]���Єy���h-�A�""t�N�$��L�$t�i��g��
O]�g�j'W�A!�Aġ���Ap��t!�x�m?��{��_a��������V����G�|g�8���y�X�'' 1�.%I���t����&!�/�>���+�'j�[�X�W��5�\�KZ��V��ۢ����o����&�s5�d�OY�__o���L[R��eݤY�3�vsp�bwհ;�P��@ǽ��!5N����w��T�)\W@�D+h"�
�+���tT�典#��1�&]��bd0�O���i95��R�L���ע�'v{+�nQ����9%2�C�hJ��=����t0E~%�S#ea��dn��;N�\SxW6�CuO�]����D�>x
�CC�-'��O�>����0EO��C �1\��_���z��d�T�@;1�2R�Э�.g3�X�ı�G>6�%�y�햗��ٔչw��%1��يC��e7��5�2*܍�5 ����}2���F�Ҍ��|��+��\Y.�8աD��e��;�ؗD���:s�m䜣�g DF����k+�4�3�1��)�����Qd:�ق�+��<���1"�5V�V���c���C���uQ�� y�$]z�6Zs�<�����h>�0��"��b��b��p>��ҩ�e�>Ι�{~�}��bO�z�<�� ��)<��^��g0�V��+N�((��3I,��q����1�8��l>��GX ���6�oL��f�$0�g���ɶJ#���N���/VK$����۫��͡y�ϛ"�g�b��S�I�2�خ
�y��ˌ��� �4�����f9u����~�E��מy0�j�߈��G����d7*w�տ�Ed���1'���_o�1���[^��s��Z�~��)��$d�$��D�3��@���Ɍꍳ�=�x(=��%WqߤO�Vw6H��_|�x�-����F��jjik�����"�N�s�\�x�4�H�/�؃X�����Sȭ�:;g,�����ԧ��	~�A���V��v; [���������U�n�"����?��wlPFf5�WF���=`�F����N؄'g��k�
�zT^֙�����'Ol�z�I���0��Г�mZmԦgd�r/ _l�&o�,t�P��_D��l�><�����m73�C��%�#���y8/V�^��*"n�EEtxx�u6r�F΂�[^ʦ@3�?��"�a�uʛ3��+(ѭlb�+c�'da�3�i���NY�]�~�p3ᇽz��:�'V��ߡg�E�!W��E(5޳e[��Q��s�`�c3�#�'��r�T|yY ���%%��N$"�&�6��4S<�Lq��U`}wSD6����~��!��Hw�ѹU>=Z�n�W���In�	Hv/�}�e��t�]j��!E���V*~��v�_�UZ�}U&N	!�ȖȠ9q��d����ҴvU��o�]F���DP���Y� ɤ��_����y�;4��4�kXo�J���$Ccg� �Y۫)��k!/�a��Wv��1���(b����ăm����!�dٺ��խXɻp)�F'S[h�t�1���JjN��o�����C�l��v����k3~�E�=r�3�/�O��3vά���:���Z��	���C�|���r%����9��4hT�~���g��53H�{]�����4���)�<!��+]V���Oc�����$䗫dxy�����������6��R"_ó��_����̕�.���_̲/ ���7v$<M���+���o�Sڌ7*R>,���,H⾒�����Uy��3@�Y�[�I�}�^�0MwB�x%��#�<7�FU���	(Gze��$K�Yў���Rtl$���"�nS��}N7�!{�p��K��E_��0-|�#F+>?�\���2�i�v�Rmp"��j��ĉ�c,�Z -̊�q�N�o�p��Z&�u�`�}.�j��D-��:{�wA��_���ꇈJ�cD3�j�z�2�g�p�$�h1��)U��w��</'��`�w��=�<���d.���ѦhH�fOP\���9��d��8ަ&]��:�0`c�{	��"��5v��ǋ��#�j�6��@�>�Q��7ʔ�	{�AY5�"�Gl9VX3�Fŵ)���H}S
��H�!@��I��ҦZѺÍ���'�f4��Γ�rs�5;�l-�a�WV������'��1n���S�3J~�=˼3e�Q�I0-p�AJW@�z�ۅ���{���P�#W `��"��(]FWBkT��v��\����
ZGjhg�b"y���t�������%\,A�O��a�R9nI)F���.Lb�q�c��VѓɩE�Z���\�P����D��RS��)PU'���N `^Rǉ+��Ӄ��ۥ̧
吔��Lo�ooۗ`�n�s��O��
e�h��&c�f�dL��4�N3ς���7G���S1���o~&O	���yt=�*�Հ�PxP��u>�K�������B���z*=�ح�5��u��݋0�k����{u�
kl���qDs�K�.�La���:+�֣s1V���t��41�Y�p7ߥ[H=we�$�.�9m��u��}��Qh��I�B�sH���9bMo��7�q�������יf�A�p�+,���=����1�=���4���u��ѓ�_g&��Ug���R�7�,D�E��C��P�fX'K����#ک�J�kk�Q�P���4��9������S�p�L�dk�uȜ�5ۋD&�\D+y�^�?�?kP�Atި<�iyhY��l���'(t\`����PЭb� ��H�2@�%�n��g��r�!�X �����yg��МD�:�go%+I�q���S��iC��#���ب�7�3��+P�3��<�`l"�f�uqjx�Ԓ;ۨ��fP��[��l�W�}�*?�n�0�ES�L�	��
���,������2�:Zլ�^i�{'s����Eg �p�|�)�����ɽ :�$�_�)"�%&⯗�g��ɥ�݄yY�@�p�C<��w���O�K��eh$ѓ:8M�7쀤��o��.Ԡ)��c�i�lQN��qYa>P���� �q�� L���:1�Н�I��;Lp��/E�cҚR�!����=K�R��N��v%By�'n�E�������2���Ce��ҤB{��5��J�`�.��)��}�~��F(�����ȿӡ�� �=��C1!H�rSz7�Nk�{����oM�ߌEK�q(Ɯòy;�˵���,�`X������z�a����9�#a�kq����w>�٬���V�����S�@�8n;�}~�bR�bt���+�@�B��8�ہ�֎m���[(x�Q��	1�7�S9� �~5Cw&-�X>�����fV��H�t��#���w�+���rn�? %��|�.�P��AԎ��Z٠�&L )�?�~`~�����!d�=|��+#~D�}}ᱍ���$%��r���#g�կ8�$"�Ma�iP(D%@�l�mG��uŊ�7�!Bn8�β�fJ��[Mr�n�t�^gu�m^�eM�/k�j}00�A�㩙�Cvm<R׫-R1QJε�A�K�M�>|K(y6C~4w6�i��Z���,���rW�`�쁤��4�u������Ck���q�^t6Bo�m��9�F�7/�N���!�d�����42��V>U��CSW�9���&peV��j�\;v�	H�}o�g�=nQ(��%��9~GE��cޞ8���U�_��\l�Ji}���@q��/L���%���?����m"tu��#6�&E3��ךY����\��Ԋ,'2�����󼘊Y�A4�:)�h���*w�}Ȧ������Ѱ㋴�4��_��i��X�^8v���� A�0���;I�n2�{.��6�Ơ3�ɢ��Jj��=�S�
8bJ�4}Ђ�I�AG�A�0�p�+�.Cy �70hyo�`\i�Y���T.��m�Ц,2�8M�?�1+���@�X�!w�~A�O���ge�=uR2���Ghc$�-O#	eľ�cdۙ9��ׅ�����yG�L@����A�j���{7 =��=U�7�)��P��8;˴Բo�d���J���n������k��[�.����5��� G�7�<������p&�Gkm��i71�	^�H��#�vGO����M��T��Q�޻J
��f-�Z)�%��dݮ�J��:��x_Wr`���j�<�6(��Z���~}���z�>�0N�$,p�Ϡ����֣̑j�a�Ħq���7r��ݭjsЋ��c��N�P���*��T��W~�n�>k�0 ��t<i�=r
zl#P^���G�tF��Z��꛳������!ZeKv%�x�����ׁ��R�iT8/,L���O
?�	�c�1m�%�C�~��T��97(����������zd�>�*��}��/dn��k�_���{[A~�q���o��*��Ⱥ�¤F���N�v�O�<sɿ�I9L tlg��HnMÀ�i�%�w'!0S��